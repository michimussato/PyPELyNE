MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       5��Aq��q��q����p��x�[��x�	��VX�r��q��$��x� K��x�p��x�p��Richq��                PE  L ۪�O        � !	  �  �      "                                                             P� M   �� (                            � p  `                            �� @                                       .text   E�     �                   `.rdata  ��     �   �             @  @.data   �3   �     �             @  �.reloc  P&   �  (   �             @  B                                                                                                                                                                                                                                                                                                                                                                                                U��`�V��H�QV�ҡ`��H�U�AVR�Ѓ���^]� U��`�V��H�QV�ҡ`��U�H�E�IRj�PV�у���^]� ����������U��`��H�A�U���R�Ћ`��Q�Jj j��E�h P�эU�R�  �`��H�A�U�R�Ћ`��Q�J�E�P�ы`��B�Pj j��M�h�Q�ҍE�P�n  �`��Q�J�E�P�у�8��  ��uP�`��B�P�M�Q�ҡ`��H�Aj j��U�h�R�ЍM�Q�  �`��B�P�M�Q�҃�3���]á`��H�A�U�R�Ћ`��Q�Jj j��E�h�P�эU�R��  �`��H�A�U�R�Ћ`��Q�J�E�P�ы`��B�Pj j��M�h Q�ҍE�P�  �`��Q�J�E�P�у�8�   ��]�����������������������U��E��P=�  SV��  t/�� t���)  �d��R  ���^��[��]�^�   [��]ËE3�9��  W�@�<� �<��[  �7�h�Ƌ��:u��t�P:Qu������u�3����������   �`�Ɗ:u��t�P:Qu������u�3����������   �X�Ɗ:u��t�P:Qu������u�3��������u3PhD�M�������M�Q�6  �`��B�P�M�Q�҃��   �4����I �:u��t�P:Qu������u�3��������uW��    �  �I�`��H�A�U�R�Ћ`��Q�Jj j��E�h P�эU�R�  �`��H�A�U�R�Ѓ��EC;�����_^3�[��]�=�  us�u��tl�~ ufj h�M��(����M�Q��$  P�U�R�E�P�O   P�9  �`��Q�J�E�P�ы`��B�P�M�Q�ҡ`��H�A�U�R�Ѓ�^3�[��]����������U��`��H�QV�uV�ҡ`��H�U�AVR�Ћ`��Q�B<�����Ћ`��Q�M�RLj�j�QP���ҋ�^]���������U��`��P�EP�EP�EP�EPQ���   �у�]� �����U���  �p�3ŉE��M�EPQ������h   R� ����|	=�  |#��`��H��0  hphH  �҃��E� �`��H�A������R�Ћ`��Q�Rj j�������P������Q�ҍ�����P��	  �`��Q�J������P�ыM�3̓����  ��]��������������U���XSVW�}���  � ��  �G$�8 ��  �G0�`��QPP�B�Ѓ�����  �M�Q�OD��z  �`��B�P4j h�  �M���h�  �M��E�   �E�    ���  �`��P�R|�E�P�M�Q�M��ҍM�舂  �`����   ��U�R�Ѓ��M�Q�OD�z  j �
  �`��B@�M�P,Q�ҋ�`��P���   ��j h�  ���Ћ`��Q�����   j h�  ���E�Ћ`��Q�����   j h�  ���E��ЋODj���j�E��y  �؉]��`��(�Q�BHj W�Ћ�����u�M���~  _^�   [��]� ��t�j���(x  �N�^�V�M�N�M�+ˍy�`��U�Q���   ����h���jBQ�E��҃��E���t��u�;u��  ���E��M�jj PWVS��w  �E�H(jWVS������E܋Ѕ���   ;]�M���   �E��������E��}��U��U��Uԅ�t4�@(�]��@0�]��@8�@X�]��E��E��]��E��E��]��E��E��]ԅ�ù} �E���E��Q�E��Qt�������ڀ}� t���Y��؀}� t���Y���M����m��n������؍M�Q�pW  �U��M���jj RWVS�*w  F;u�������E�P�GW  ���M��,}  _^3�[��]� �U��`��H�A�� �U�VR�Ћ`��Q�Jj j��E�h�P�ы`��B�P�M�Q�ҡ`��H�Aj j��U�h�R��j j j �M�Qh� j �U�RhЫ ��  ��`��H�A�U���HR�Ћ`��Q�J�E�P�у���^��]ø   � ��������U��V���UP  �Et	V�Y  ����^]� ���������������Vh�jh��j�,Z  ������t����O  ���^�3�^���������������U��E�`�� ]��U��`��P8�EPQ�JD�у�]� ���̡`��H8�Q<�����U��`��H8�A@V�u�R�Ѓ��    ^]�������������̡`��H8�������U��`��H8�AV�u�R�Ѓ��    ^]��������������U��`��P8�EP�EP�EPQ�J�у�]� ������������U��`��P8�EP�EPQ�J�у�]� �`��P8�BQ�Ѓ����������������U��`��P8�EPQ�J �у�]� ����U��`��P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U��`��P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U��`��P8�EP�EPQ�J(�у�]� U��`��P8�EP�EP�EPQ�J,�у�]� ������������U��`��P8�EP�EP�EPQ�J�у�]� ������������U��`��P8�EP�EP�EP�EP�EPQ�J�у�]� ����U��`��P8�EP�EPQ�J0�у�]� U��`��P8�EP�EP�EPQ�J4�у�]� ������������U��`��P8�EPQ�J8�у�]� ����U��`��H��x  ]��������������U��`��H��|  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H�A,]�����������������U��`��H���  ]��������������U��`��H�QV�uV�ҡ`��H�Q8V�҃���^]�����̡`��H�Q<�����U��`��H�I@]����������������̡`��H�QD����̡`��H�QH�����U��`��H�AL]�����������������U��`��H�IP]�����������������U��`��H��<  ]��������������U��`��H��,  ]��������������U��`��H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡`��H���   ��`��H���  ��U��`��H�U�ER�UP�ER�UP���   Rh�2  �Ѓ�]����������������U��`��H�A]�����������������U��`��H��\  ]��������������U��`��H�AT]�����������������U��`��H�AX]�����������������U��`��H�A\]����������������̡`��H�Q`�����U��`��H���  ]�������������̡`��H�Qd����̡`��H�Qh�����U��`��H�Al]�����������������U��`��H�Ap]�����������������U��`��H�At]�����������������U��`��H��D  ]��������������U��`��H��  ]��������������U��`��H�Ix]�����������������U��`��H��@  ]��������������U��V�u���B  �`��H�U�A|VR�Ѓ���^]���������U��`��H���   ]��������������U��`��H��h  ]��������������U��`��H��d  ]��������������U��`��H���  ]�������������̡`��H���   ��U��`��H��l  ]��������������U��`��H��   ]��������������U��`��H��  ]��������������U��V�u���Rs  �`��H���   V�҃���^]���������̡`��H��`  ��U��`��H��  ]��������������U��`��H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U��`��H���  ]��������������U��U�E�`��H�E���   R���\$�E�$P�у�]�U��`��H���   ]��������������U��`��H���   ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���   ]��������������U��`��H���   ]��������������U��`��H���   ]��������������U��`��H���   ]��������������U��`��H���   ]��������������U��`��H���   ]��������������U��`��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��`��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��`��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��`��H��8  ]��������������U��V�u(V�u$�E�@�`��R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@�`��R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��`��P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U��`��P0�EP�EP�EP�EPQ���   �у�]� ����̡`��P0���   Q�Ѓ�������������U��`��P0�EP�EPQ���   �у�]� �������������U��`��P0�EP�EP�EP�EPQ���   �у�]� ����̡`��P0���   Q�Ѓ������������̡`��H0���   ��U��`��H0���   V�u�R�Ѓ��    ^]�����������U��`��H��H  ]��������������U��`��H��T  ]�������������̡`��H��p  ��`��H���  ��U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �`����   �Qj PV�ҡ`����   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M���l  P�E�hicMCP�k������M���l  �`����   �JT�E�P�у���u(�u���jl  �`����   ��M�Q�҃���^��]á`����   �AT�U�R�Ћu��P���jl  �`����   �
�E�P�у���^��]�������������U��`��H��  ]��������������U��`��H��\  ]��������������U��`��H�U��t  ��V�uVR�E�P�у����  �M��K  ��^��]�����U��`��H�U���  ��VWR�E�P�ы`��u���B�HV�ы`��B�HVW�ы`��B�P�M�Q�҃�_��^��]����������������U��`��H�U���  ��VWR�E�P�ы`��u���B�HV�ы`��B�HVW�ы`��B�P�M�Q�҃�_��^��]����������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H�U�E��VWj R�UP�ERP��t  �U�R�Ћ`��Q�u���BV�Ћ`��Q�BVW�Ћ`��Q�J�E�P�у�(_��^��]��U��`��H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �`����   j P�BV�Ћ`����   �
�E�P�у�$��^��]���U��`��H��8  ]��������������U���  �p�3ŉE��M�EPQ������h   R���  ����|	=�  |#��`��H��0  hphH  �҃��E� �`��H��4  ������Rh��ЋM�3̓���  ��]�������U��`��H��  ��V�U�WR�Ћ`��Q�u���BV�Ћ`��Q�BVW�Ћ`��Q�J�E�P�у�_��^��]����U��`��H��  ��V�U�WR�Ћ`��Q�u���BV�Ћ`��Q�BVW�Ћ`��Q�J�E�P�у�_��^��]����U��`��H��p  ��$�҅�trh���M��g  �`��P�E�R4Ph���M��ҡ`��P�E�R4Ph���M���j �E�P�M�hicMCQ�����`����   ��M�Q�҃��M��g  ��]�U��`��H��p  ��$V�҅�u�`��H�u�QV�҃���^��]�Wh!���M���f  �`��P�E�R4Ph!���M���j �E�P�M�hicMCQ�����`����   �QHP�ҋu���`��H�QV�ҡ`��H�QVW�ҡ`����   ��U�R�Ѓ�$�M��f  _��^��]������U��`��H��p  ��$V�҅�u�`��H�u�QV�҃���^��]�Wh����M��,f  �`��P�E�R4Ph����M���j �E�P�M�hicMCQ�����`����   �QHP�ҋu���`��H�QV�ҡ`��H�QVW�ҡ`����   ��U�R�Ѓ�$�M���e  _��^��]������U��`��H��p  ��$�҅�u��]�Vh#���M��te  �`��P�E�R4Ph#���M���j �E�P�M�hicMCQ������`����   �Q8P�ҋ�`����   ��U�R�Ѓ��M��Ue  ��^��]���������������U��`��H��p  ��$�҅�u��]�Vhs���M���d  �`��P�E�R4Phs���M���j �E�P�M�hicMCQ�W����`����   �Q8P�ҋ�`����   ��U�R�Ѓ��M��d  ��^��]���������������U��`��H���  ]��������������U��`��H��@  ]��������������U��`��H���  ]��������������U��V�u���t�`��QP��D  �Ѓ��    ^]������U��`��H��H  ]��������������U��`��H��L  ]��������������U��`��H��P  ]��������������U��`��H��T  ]��������������U��`��H��X  ]��������������U��`��H��\  ]�������������̡`��H��d  ��U��`��H��h  ]��������������U��`��H��l  ]�������������̡`��H���  ��U��`��H�U���  ��VR�E�P�ыu��P���b  �M��b  ��^��]�����U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H��l  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H��$  ]��������������U��`��H��(  ]��������������U��`��H��,  ]�������������̡`��H��0  ��`��H��<  ��U��`��H���  ]�������������̡`��H���  ��U��`��H���  ]������������������������������U��`��H��  ]�������������̡`��H��P  ��U��`��H��`  ]�������������̡`����   ���   ��Q��Y��������U��`��H�A�U��� R�Ћ`��Q�Jj j��E�h�P�ыUR�E�P�M�Q�]����`��B�P�M�Q�ҡ`��H�A�U�R�Ћ`��Q�J�E�P�у�,��]��U��`��P�EP�EP�EPQ�J�у�]� �����������̡`�V��H�QV�ҡ`��H$�QDV�҃���^�����������U��`�V��H�QV�ҡ`��H$�QDV�ҡ`��U�H$�AdRV�Ѓ���^]� ��U��`�V��H�QV�ҡ`��H$�QDV�ҡ`��U�H$�ARV�Ѓ���^]� ��U��`�V��H�QV�ҡ`��H$�QDV�ҡ`��H$�U�ALVR�Ѓ���^]� �̡`�V��H$�QHV�ҡ`��H�QV�҃�^�������������U��`��P$�EPQ�JL�у�]� ����U��`��P$�R]�����������������U��`��P$�Rl]����������������̡`��P$�Bp����̡`��P$�BQ�Ѓ����������������U��`��P$��VWQ�J�E�P�ы`��u���B�HV�ы`��B�HVW�ы`��B�P�M�Q�҃�_��^��]� ���U��`��P$�EPQ�J�у�]� ����U��`��P$��VWQ�J �E�P�ы`��u���B�HV�ы`��B$�HDV�ы`��B$�HLVW�ы`��B$�PH�M�Q�ҡ`��H�A�U�R�Ѓ� _��^��]� ���U��`��P$��VWQ�J$�E�P�ы`��u���B�HV�ы`��B$�HDV�ы`��B$�HLVW�ы`��B$�PH�M�Q�ҡ`��H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e����`��Q$�JH�E�P�ы`��B�P�M�Q�҃���^��]� ����̡`��P$�B(Q��Yá`��P$�BhQ��Y�U��`��P$�EPQ�J,�у�]� ����U��`��P$�EPQ�J0�у�]� ����U��`��P$�EPQ�J4�у�]� ����U��`��P$�EPQ�J8�у�]� ����U��`��UV��H$�ALVR�Ѓ���^]� ��������������U��`��H�QV�uV�ҡ`��H$�QDV�ҡ`��H$�U�ALVR�Ћ`��E�Q$�J@PV�у���^]�U��`��UV��H$�A@RV�Ѓ���^]� ��������������U��`��P$�EPQ�J<�у�]� ����U��`��P$�EPQ�J<�у����@]� ���������������U��`��P$�EP�EPQ�JP�у�]� U��`��P$�EPQ�JT�у�]� ���̡`��H$�QX�����U��`��H$�A\]�����������������U��`��P$�EP�EP�EPQ�J`�у�]� �����������̡`��H(�������U��`��H(�AV�u�R�Ѓ��    ^]��������������U��`��P(�R]����������������̡`��P(�B�����U��`��P(�R]�����������������U��`��P(�R]�����������������U��`��P(�R ]�����������������U��`��P(�E�RjP�EP��]� ��U��`��P(�E�R$P�EP�EP��]� �`��P(�B(����̡`��P(�B,����̡`��P(�B0�����U��`��P(�R4]�����������������U��`��P(�RX]�����������������U��`��P(�R\]�����������������U��`��P(�R`]�����������������U��`��P(�Rd]�����������������U��`��P(�Rh]�����������������U��`��P(�Rl]�����������������U��`��P(�Rx]�����������������U��`��P(���   ]��������������U��`��P(�Rt]�����������������U��`��P(�Rp]�����������������U��`��P(�BpVW�}W���Ѕ�t:�`��Q(�Rp�GP���҅�t"�`��P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U��`��P(�BtVW�}W���Ѕ�t:�`��Q(�Rt�GP���҅�t"�`��P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U����`��E�    �E�    �P(�RhV�E�P���҅���   �E���uG�`��H�A�U�R�Ћ`��Q�E�RP�M�Q�ҡ`��H�A�U�R�Ѓ��   ^��]� �`��Qh�he  P���   �Ћ`����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P��.  ��3�^��]� �M��U�j IQ�MR������E�P�.  ���   ^��]� ���������������U��`���V��H�A�U�R�Ѓ��M�Q������^��u�`��B�P�M�Q�҃�3���]� �`��H$�E�I�U�RP�ы`��B�P�M�Q�҃��   ��]� �U��Q�`��P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U��`��P(�R8]�����������������U��`��P(�R<]�����������������U��`��P(�R@]�����������������U��`��P(�RD]�����������������U��`��P(�RH]�����������������U��`��P(�E�R|P�EP��]� ����U��`��P(�RL]�����������������U��`��E�P(�BT���$��]� ���U��`��E�P(�BPQ�$��]� ����̡`��H(�Q�����U��`��H(�AV�u�R�Ѓ��    ^]��������������U��`��P(���   ]��������������U��`��H(�A]����������������̡`��H,�Q,����̡`��P,�B4�����U��`��H,�A0V�u�R�Ѓ��    ^]�������������̡`��P,�B8�����U��`��P,�R<��VW�E�P�ҋu���`��H�QV�ҡ`��H$�QDV�ҡ`��H$�QLVW�ҡ`��H$�AH�U�R�Ћ`��Q�J�E�P�у�_��^��]� �������U��`��P,�E�R@��VWP�E�P�ҋu���`��H�QV�ҡ`��H�QVW�ҡ`��H�A�U�R�Ѓ�_��^��]� ��̡`��H,�j j �҃��������������U��`��P,�EP�EPQ�J�у�]� U��`��H,�AV�u�R�Ѓ��    ^]�������������̡`��P,�B����̡`��P,�B����̡`��P,�B����̡`��P,�B ����̡`��P,�B$����̡`��P,�B(�����U��`��P,�R]�����������������U��`��P,�R��VW�E�P�ҋu���`��H�QV�ҡ`��H$�QDV�ҡ`��H$�QLVW�ҡ`��H$�AH�U�R�Ћ`��Q�J�E�P�у�_��^��]� �������U��`��H��D  ]��������������U��`��H��H  ]��������������U��`��H��L  ]��������������U��`��H�I]�����������������U��`��H�A]�����������������U��`��H�I]�����������������U��`��H�A]�����������������U��`��H�I]�����������������U��`��H���  ]��������������U��`��H�A]�����������������U���V�u�E�P��������`��Q$�J�E�P�у���u-�`��B$�PH�M�Q�ҡ`��H�A�U�R�Ѓ�3�^��]Ë`��Q�J�E�jP�у���u=�U�R��������u-�`��H$�AH�U�R�Ћ`��Q�J�E�P�у�3�^��]Ë`��B�HjV�у���u�`��B�HV�у����I����`��Q$�JH�E�P�ы`��B�P�M�Q�҃��   ^��]�����������U��`��H�A ]�����������������U��`��H�I(]�����������������U��`��H��  ]��������������U��`��H��   ]��������������U��`��H��  ]��������������U��`��H��  ]��������������U��`��H�A$��V�U�WR�Ћ`��Q�u���BV�Ћ`��Q$�BDV�Ћ`��Q$�BLVW�Ћ`��Q$�JH�E�P�ы`��B�P�M�Q�҃�_��^��]������U��`��H���  ��V�U�WR�Ћ`��Q�u���BV�Ћ`��Q$�BDV�Ћ`��Q$�BLVW�Ћ`��Q$�JH�E�P�ы`��B�P�M�Q�҃�_��^��]���U��`��H���  ]��������������U���<���SVW�E�    ��t�E�P�   �������/�`��Q�J�E�P�   �ы`��B$�PD�M�Q�҃��}�`��H�u�QV�ҡ`��H$�QDV�ҡ`��H$�QLVW�҃���t)�`��H$�AH�U�R����Ћ`��Q�J�E�P�у���t&�`��B$�PH�M�Q�ҡ`��H�A�U�R�Ѓ�_��^[��]���U��`��H�U���  ��VWR�E�P�ы`��u���B�HV�ы`��B$�HDV�ы`��B$�HLVW�ы`��B$�PH�M�Q�ҡ`��H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]��������������U��`��H���  ]�������������̡`��H���   ��U��`��H���   V�uV�҃��    ^]�������������U��`��P�]��`��P�B����̡`��P���   ��U��`��P�R`]�����������������U��`��P�Rd]�����������������U��`��P�Rh]�����������������U��`��P�Rl]�����������������U��`��P�Rp]�����������������U��`��P�Rt]�����������������U��`��P���   ]��������������U��`��P��  ]��������������U��`��P�Rx]�����������������U��`��P���   ]��������������U��`��P�R|]�����������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P�EPQ��  �у�]� �U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��E��t �`��R P�B$Q�Ѓ���t	�   ]� 3�]� U��`��P �E�RLQ�MPQ�҃�]� U��E��u]� �`��R P�B(Q�Ѓ��   ]� ������U��`��P�R]�����������������U��`��P�R]�����������������U��`��P�R]�����������������U��`��P�R]�����������������U��`��P�R]�����������������U��`��P�R]�����������������U��`��P�E�R\P�EP��]� ����U��`��P�E��  P�EP��]� �U��`��E�P�B ���$��]� ���U��`��E�P�B$Q�$��]� �����U��`��E�P�B(���$��]� ���U��`��P�R,]�����������������U��`��P�R0]�����������������U��`��P�R4]�����������������U��`��P�R8]�����������������U��`��P�R<]�����������������U��`��P�R@]�����������������U��`��P�RD]�����������������U��`��P�RH]�����������������U��`��P�RL]�����������������U��`��P�RP]�����������������U��`��P���   ]��������������U��`��P�RT]�����������������U��`��P�EPQ��  �у�]� �U��`��P���   ]��������������U��`��P���   ]��������������U��`��P�RX]����������������̡`��P���   ��U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]��������������U��`��P���   ]�������������̡`��P���   ��U��`��P���   ]�������������̡`��P���   ��`��P���   ��`��P���   ��U��`��H���   ]��������������U��`��H��   ]��������������U��`��H�U�E��VWRP���  �U�R�Ћ`��Q�u���BV�Ћ`��Q�BVW�Ћ`��Q�J�E�P�у�_��^��]������������U��`��H���  ]��������������U��`��P(�BPVW�}�Q�]���E�$�Ѕ�tM�`��G�Q(�]�E�BPQ���$�Ѕ�t,�`��G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U��`��P(�BTVW�}����$���Ѕ�tE�`��G�Q(�BT�����$�Ѕ�t(�`��G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U��`��P(�} �R8����P��]� �U��`��P�BdS�]VW��j ���Ћ`��Q�����   h�Fh�  V�Ћ`����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ`��Q(�BHV���Ѕ�t �`��Q(�E�R VP���҅�t�   �3��EP�  ��_��^[]� ������U���V�E���MP�k���P���#����`��Q�J���E�P�у���^��]� ���U��`��P�E���   ��VWP�EP�E�P�ҋu���`��H�QV�ҡ`��H�QVW�ҡ`��H�A�U�R�Ѓ�_��^��]� ������������U��E��u�d��MP�EPQ�#?  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3hj;h��j�]  ����t
W���^����3��F��u_^]� �~ t3�9_��^]� �`��H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   �`��H<�Q��3Ʌ����^��������������̃y t�   ËA��uË`��R<P��JP�у��������U����u�`��H�]� �`��J<�URP�A�Ѓ�]� ���������������U��d���u�`��H�]Ë`��J<�URP�A�Ѓ�]�U��d���$V��u�`��H�1��`��J<�URP�A�Ѓ����`��Q�J�E�SP�ы`��B�P�M�QV�ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@�� j �M�Q�U�R�M��Ћ`��Q�J���E�P���у���[t.�`��B�u�HV�ы`��B�P�M�Q�҃���^��]á`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�u�QV�ҡ`��H�A�U�VR�Ћ`��Q�J�E�P�у���^��]���������������U��d���$SV��u�`��H�1��`��J<�URP�A�Ѓ����`��Q�J�E�P�ы`��B�P�M�QV�ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@�� j �M�Q�U�R�M��Ћ`��Q�J���E�P���у���t/�`��B�u�HV�ы`��B�P�M�Q�҃���^[��]á`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@��j �M�Q�U�R�M��Ћ`��Q�J���E�P���у����3����`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�u�QV�ҡ`��H�A�U�VR�Ћ`��Q�J�E�P�у���^[��]����������������U��d���$SV��u�`��H�1��`��J<�URP�A�Ѓ����`��Q�J�E�P�ы`��B�P�M�QV�ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@�� j �M�Q�U�R�M��Ћ`��Q�J���E�P���у���t/�`��B�u�HV�ы`��B�P�M�Q�҃���^[��]á`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@��j �M�Q�U�R�M��Ћ`��Q�J���E�P���у����3����`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@��j �M�Q�U�R�M��Ћ`��Q�J���E�P���у���������`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҋu�E�P���#����`��Q�J�E�P�у���^[��]�������U��d���$SV��u�`��H�1��`��J<�URP�A�Ѓ����`��Q�J�E�P�ы`��B�P�M�QV�ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@�� j �M�Q�U�R�M��Ћ`��Q�J���E�P���у���t/�`��B�u�HV�ы`��B�P�M�Q�҃���^[��]á`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@��j �M�Q�U�R�M��Ћ`��Q�J���E�P���у����3����`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M��ҡ`��H�A�U�R�Ћ`��Q�Jj j��E�h\P�ы`��B�@@��j �M�Q�U�R�M��Ћ`��Q�J���E�P���у���������`��P�E��RHjP�M��ҡ`��P�E�M��RLj�j�PQ�M���j h\�M��¬���`��P�R@j �E�P�M�Q�M��҅��`��H�A�U�R���Ѓ���t/�`��Q�u�BV�Ћ`��Q�J�E�P�у���^[��]Ë`��M��B�PHjQ�M��ҡ`��P�E�M��RLj�j�PQ�M��ҋu�E�P�������`��Q�J�E�P�у���^[��]���������������U��`��H<�A]����������������̡`��H<�Q�����V��~ u>���t�`��Q<P�B�Ѓ��    W�~��t�������W�  ���F    _^��������U���V�E�P���������P��������M��������^��]��̃=l� uK�d���t�`��Q<P�B�Ѓ��d�    �p���tV���@���V�*  ���p�    ^������������U���8�`��H�AS�U�V3�R�]��Ћ`��Q�JSj��E�h`P�ы`��B<�P�M�Q�ҋ�`��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��J  �M�Q�U�R�M��K  ����   W�}�}���   �`����   �U��ATR�Ћ�����tB�`��Q�J�E�P���у��U�Rj�E�P�������`��Q�ȋBxW���E���t�E� ��t�`��Q�J�E�P����у���t�`��B�P�M�Q����҃��}� u"�E�P�M�Q�M��?J  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_�`��H�A�U�R�Ћ`��Q�JSj��E�h`P�ы`��B<�P�M�Q�ҋ�`��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��1I  �M�Q�U�R�M��I  ���p  W�}��I �E����   �`����   �U��ATR�Ћ�������   �`��Q�J�E�P���ы`��B���   ���M�Qj�U�R���Ћ`��Q�J���E�P�ы`��B�P�M�QV�ҡ`��H�A�U�R�Ћ`��Q�Bx��W�M����E��t�E ��t�`��Q�J�E�P����у���t�`��B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�`����   P�BH�Ћ`��Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��"H  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��G  �EP�M�Q�M�u��u��G  ����   �u���E���tA��t<��uZ�`����   �M�PHQ�ҋ`��Q���ȋBxV�Ѕ�u-�   ^��]Ë`����   �E�JTP��VP�[�������uӍUR�E�P�M��DG  ��u�3�^��]����������V��~ u>���t�`��Q<P�B�Ѓ��    W�~��t������W�t	  ���F    _^�������̋�� p���������p���������̅�t��j�����̡`��P��  ��`��P��(  ��U��`��P��   ��V�E�P�ҋuP�������M��������^��]� ��������̡`��P��$  ��U��`��H��  ]��������������U��`��H���  ]�������������̡`��H��  ��U��`��H���  ]��������������U��`��H��x  ]��������������U��`��H��|  ]�������������̡`��H��d  ��U��`��H��p  ]��������������U��`��H��t  ]��������������U���EV���pt	V�  ����^]� �������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���D  �����   �ESP�M�������`��Q�J�E�P�ы`��B�Pj j��M�htQ�҃��E�P�M�����j j��M�Q�U�R��d���P������P�M�Q�w�����P�U�R�j������P��E  ���M���������M��������d���������M�������`��H�A�U�R�Ѓ��M�������[t	V��C  ����^��]� ���U��EVP���N  �����^]� �����Q�C  Y���������U��E�M�U�H4�M�P �U��M�@ j �@8po �@<�o �@@�o �@D0o �@H�o �@L�o �@P@o �@l�o �@Xp �@\Po �@`�o �@d�o �@T p �@h�o �@p o �@t`o �P0�H(�@,    ]��������������U���   h�   ��`���j P�ē  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj������8��]��������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U��V�u���t�`��QP��Ѓ��    ^]���������̡`��H��@  hﾭ���Y����������U��E��t�`��QP��@  �Ѓ�]����������������U��`��H���  ]��������������U��`��H��  ]�������������̡`��H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�1�  ������u_^]Ã} tWj V�L�  ��_������F�t�   ^]���U��`��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW赑  ������u_^]�Wj V�֐  ��_������F�t�   ^]�������������U��`��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�5�  ������u_^]�Wj V�V�  ��_������F�t�   ^]�������������U��`��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW赐  ������u_^]�Wj V�֏  ��_������F�t�   ^]�������������U��`��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�5�  ������u_^]�Wj V�V�  ��_������F�t�   ^]�������������U��M��t-�=t� t�y���A�uP衐  ��]á`��P�Q�Ѓ�]��������U��M��t-�=t� t�y���A�uP�a�  ��]á`��P�Q�Ѓ�]��������U��`��H�U�R�Ѓ�]���������U��`��H�U�R�Ѓ�]���������U��`��E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��  ������u_^]�Wj V��  ��_������F�t�   ^]���������U��`��E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   �`���t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��  ������u_^]�Wj V�#�  ��_������F�t�   ^]����������U��E��w�   �`���t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�o�  ������u_^]�Wj V萌  ��_������F�t�   ^]�������U��`��H�U�R�Ѓ�]���������U��`��H�U�R�Ѓ�]���������U��`��H�U�R�Ѓ�]���������U��`��H�U�R�Ѓ�]���������U�����E��������u
����]���������u
���x]�]��  ����U��V�u�F��F����������������茒  ����������D�Ez��^��P�X]��������������N�X�N^�X]��������P�P�P�P �P(�P0�P8�P@�PH�PP�PX����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U�������M�P�P�P�P �P(�P0�P8�P@�PH�PP�XX���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��V�u�������E���P�V�H�N�P�V�H�N�P�V��^]���������U��V�u���r����E� �^�@�^8�@���^X^]����������U���V�u���?����E�'�  �]��E��  �E��VX�������^@���^P�^8^��]�U���V�u��������E��  �]��E謋  �E��V�������^H���^(�^X^��]�U���V�u�������E觌  �]��E�l�  �E��V�����V0���^ �^8^��]���U�������e�5��U��$聐  �m����������E���������Az
���.���]��؋�]��������������U���`�E��P�MЋH�M؋H�UԋP�M��M�U܋P�U��w=�$��{ � �����@�����`���]��6����� �@���@�����]��� �������`�@�����]����]�VW�}�]�����u��$������]��G�u��$������]��u��G�$������]ȍu���$������]��u��G�$�����]��u��G�$�����E�����_�E�^�����������E����E������E�����������A�Eu�E���E��X�E��X��]ËMЋUԉ�M؉P�U܉H�M��P�U�H�P��]ÍI fz Kz �z fz Kz �z ��������U�����V�u��VW�}�^�G����������ƍ  �U���������Au>�����W��������z��_����^�^^��]��x_����^�^^��]�����_���?�$��z	�m�������d���������G�u���  �^��_�^��^��]���������������U���hV�u�FP�M�Q�Y����V0R�E�P�L�����H�M�VQ�?����E��^���A  �$�� �E������$��������U��]�  ����������Au�E��E��;�  �]��E��  ���]��E��E�� �  ���]�����z�-��E��  �E����$�n������U���  ��������Au%�E����E��ѐ  �]��E����E����  �E��c  ���]��E����E���襐  ���]�����Au��-��E��5  �E������$��������U��v�  ��������Au0�E��E��V�  �]��E��E��H�  �E�E����X�E��X��]����]��E����E���  ���]�����Au���E�E����X�E��X��]��EЃ����$�`������U���  ����������Au0�E��E��Ï  �]��E��E�赏  �E�E����X�E��X��]����]��E��E�莏  ���]������m������E�E�����X�E��X��]��E؃��$��������U��N�  ��������Au4�E����E��,�  �]��E����E���  �E�E����X�E��X��]����]��E����E�����  ���]�����A������%��E�E�����X�E��X��]��E����$�,������U�豆  ��������Au:�E����E�菎  �]��E����E���  �]��E��E�E�����X�E��X��]����]��E��E��R�  ���]�����A�4������E���  �E����E�����草  �U���������A��   �������U��E����E��E���������������Az�����.��������u
�����������訌  �E��E������U����U�����z'�����������<  �������]��,  �x��������A�  �������]��  ����]����}��$��z	��������������U�����������Au���]�����E��u��?�  �]��E���  �]��E��Ƀ  �E��M��E������������M�����������Az�����$��������u
�������萋  �����U����]�����z#�-��E�]��E��E�����X�E��X��]ËE���E��E�����X�E��X��]��ڋE������X�E��X��]Ë��| $} �} f 0~ �~ ������������U�����   V���u�����Dz%�V����Dz�^����Dz�u���������^��]����W�}�U�衂  ��u)�]��E����  �]��F�U�胂  �]��E�訃  �]��'�]��E�蘃  �]��F�U��Z�  �]��E���  �]��F�U��A�  �]��E��f�  ����  �$�\� �E��u���E��E�P�ɍM��E�Q�ˍU�R��p�����P�E��������������]������������]��E������]������]������]��E����]������������]��������������]����]���ݕp���ݕx����]��9���_��^��]��E���p�����Q�E؍U���R�E�E���P�ˍM�Q�U�������ݝp����E����E���������ݝx��������E������]��E��]������]��������]��������]������������]��+  ����p����E�R�ɍE��E�P���M���Q�U�R�U�����ݝp����E����E�����ݝx����E������]������]������������]��E����������]������]������������]����  �E���p�����P�E��M���Q�E��U���R�ˍE�P�U��E������E�������ݝp�������ݝx����E����������]������������]��������]������������]����]��E����]����   �E���p�����Q�E�U���R�E��E���P�ʍM��E�Q����������ݝp�������������ݝx������E������]������������]������������]��������]������]������]��E��   ����p����E�R�ɍE��E�P���M���Q�U�R�]��E����E�������ݝp�����ݝx������E������]������������]������]��������������]������E����������]��������]������������u�]�����U��U��]��^���_��^��]Ë�ڂ � � �� �� � ������������U���xV�uW�   �}��E��P�M�Q�>�����H�U��P�M��H�U��P�@�M��M��U�Q�U�R�E�������P�M��H�U��P�M��H�UċP�EЉM�P�M�Q�U�������E���E��H�UЋP�MԋH�U؋P�@�E�U��E������M�������������u�������������u
�����褅  �}�u��EȍM��e�VQ��E��e��^�E��e��^�H�������H�N�P�V�H�N�P�V�@�F�������Dz,�V����Dz"�V����Dz����������^�^�_^��]�_��^��]�����U���0V�uW���.�����}�������Dz�W����Dz
�W����D{�E��������Dz
_�؋�^��]����U��|  �]��E���}  �]��E�WP�l���� �E������@���@�������������������E������]������]������������]��������������������������]��E����]����E������]��E��^�E��^ �E��^(�E������]��������������]����E�����_�]����E��^0�E��^8�E��^@���������������^H���^P�^X^��]��������������U��E�A    �]� �������������U��Q�@i�� %����E���E���}���5���]���U��Q�@i�� %����E���E���}���5����%���]�����������U���V��~ ��   �����������؍Ai�� %����ȉM��E���}����Hi�� ���������U��щU��E���}���������U����������U�������t���������D{��ډ��������}  ���u���~  �E����F   �^^�M�������]��F�F    ��^����]�����������U���V��~ ��   �����������؍Ai�� %����ȉM��E���}����Hi�� ���������U��щU��E���}���������U����������U�������t���������D{��ډ��������|  ���u���}  �E����F   �^^�M�����]��F�F    ��^��]�������U��E�M�@�I�����A�H����� ���@�����H�E�������A�����X�i�X]�������U��E� �@�@����������Au��������������Au����������������z��������������z����������������   ��������� ������Au�E������������X�X]�������������Dz
���������5��������Dz������������������������������������5���������z���E����X�X]ËE������������P�X]�U����E� �@�U��@�U�� ��������Au�E������������X�X��]�����������Dz���������U��$�|  �E����������E����E����������������������������W�  H��wE�$�8� �����ʋE��������X�X��]��������������ۋE��������X�X��]������� � � � � ����U��M�A��A��������������������������Dz�E����P�X]ËU�؋E�� �B�`�B�`������I���I����������I���I� �����@�@�E���������j�X�j�X]�������̡`��H���   ��U��`��H���   V�u�R�Ѓ��    ^]����������̡`��H���   ��U��`��H���   V�u�R�Ѓ��    ^]����������̡`��P���   Q��Y��������������U��`��P�EPQ���   �у�]� �U��`��P�EP�EP�EP�EP�EP�EPQ���   �у�]� �������������U��`��P�EP�EP�EP�EP�EP�EPQ���   �у�]� �������������U��`��P�EP�EP�EP�EPQ���   �у�]� �����U��`��P�EP�EP�EP�EPQ��  �у�]� �����U��`��P�EP�EP�EP�EPQ���  �у�]� �����U��`��P�EP�EPQ���   �у�]� �������������U��V�uW�����  �`��H���   VW�҃�_��^]� ��U��`��P�EPQ���   �у�]� �U��`��P�EPQ��  �у�]� ̡`��P��0  Q�Ѓ�������������U��`��P�EP�EPQ��t  �у�]� �������������U��`��H�U���  j R�Ѓ�]���U��`��H���  V�u�R�Ѓ��    ^]�����������U��`��H���   ]��������������U��`��H���   V�u�R�Ѓ��    ^]�����������U��� ��`�3��U�Q�U�Q�]�Q�M��M��P�E�PQ�E�P�EPPP�EP�EP�EP�EPQ��d  �у�8��]��������������U��U��tA���    t8��  �M;A}*V�1�0^t	�E�    �	��  �t	�E�    ]����U��`��H��P  ]��������������U��`��H��T  ]��������������U��`��H��X  ]�������������̋��     ��������V����t�`��QP��<  �Ѓ��    ^�����������U����t�`��Q�M���  Q�MQP�҃�]� ������U����t�`��Q�M���  Q�MQP�҃�]� �����̋A@��t�`��QP�BD�Ѓ�ø   �U��`���S3�V��W�}��~D�^<�^8�^@�^H�FL   �^P�^T;���   �U�R����9  P�N�/����M��������� ;  �F�E�P����C  ��N�P�V�H�N�P�V�`��H@�Q,W�ҋ���;�tG�`��P���   Sh6  ���ЉFP�`��Q���   Sh5  ����_�FT^[��]� �F   _^[��]� ���̋��@    � d   �V����t�`��QP��<  �Ѓ��    ^�����������U��V����t�`��QP��<  �Ѓ��    �`��Q�E�MP�EQ��8  P��3҃����^��]� ��������̡`��P�BVj j����Ћ�^���������U��`��P�E�RVj P���ҋ�^]� U��`��P�E�RVPj����ҋ�^]� �`��P�B�����U��`��P���   Vj ��Mj V�Ћ�^]� �����������U��`��P�EPQ�J�у�]� ����U��`��P�EPQ�J�у����@]� ���������������U��`��P�E�RtP�ҋ`����   P�BX�Ѓ�]� ���U��`��P�E�Rlh#  P�EP��]� ���������������U��`��P�E�RlhF  P�EP��]� ���������������U��`��P�E�RtP�ҋ`����   �M�R`QP�҃�]� ���������������U��`��P���   ]��������������U��`��P�E���   P�҅�u]� �`����   P�B�Ѓ�]� ��������h��PhD �PN  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h��jhD �|M  ����t
�@��t]��3�]��������Vh��j\hD ���LM  ����t�@\��tV�Ѓ���^�����Vh��j`hD ���M  ����t�@`��tV�Ѓ�^�������U��Vh��jdhD ����L  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh��jhhD ���L  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh��jlhD ���lL  ����t�@l��tV�Ѓ�^�������U��Vh��h�   hD ���6L  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh��h�   hD ����K  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh��jphD ���K  ����t�@p��t�MQV�Ѓ�^]� ���^]� ��U��Vh��jxhD ���YK  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh��j|hD ���K  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh��j|hD ����J  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vh��h�   hD ���J  ����t=���   ��t3�MQ�U�VR��h��j`hD �VJ  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������h��jhD �J  ����t	�@��t��3��������������U��V�u�> t+h��jhD ��I  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h��jhD �I  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh��jhD ���II  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh��jhD ���	I  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh��j hD ����H  ����t�@ ��tV�Ѓ�^�3�^���Vh��j$hD ���H  ����t�@$��tV�Ѓ�^�3�^���U��Vh��j(hD ���iH  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh��j,hD ���H  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh��j(hD ����G  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh��j4hD ���G  ����t�@4��tV�Ѓ�^�3�^���U��Vh��j8hD ���YG  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh��j<hD ���	G  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh��jDhD ����F  ����t�@D��tV�Ѓ�^�3�^���U��Vh��jHhD ���F  ����t�M�PHQV�҃�^]� U��Vh��jLhD ���iF  ����u^]� �M�PLQV�҃�^]� �����������U��Vh��jPhD ���)F  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh��jThD ����E  ����u^Ë@TV�Ѓ�^���������U��Vh��jXhD ���E  ����t�M�PXQV�҃�^]� U��Vh��h�   hD ���E  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh��h�   hD ���6E  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh��h�   hD ����D  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���D  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���fD  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���&D  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh��h�   hD ��C  ����u�`��H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ`��Q�u���BV�Ћ`��Q�BVW�Ћ`��Q�J�E�P�у�_��^��]��U��Vh��h�   hD ���VC  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   hD ���C  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   hD ����B  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   hD ���B  ����t���   ��t�MQ����^]� 3�^]� �Vh��h�   hD ���IB  ����t���   ��t��^��3�^����������������U��Vh��h�   hD ���B  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   hD ���A  ����t���   ��t�MQ����^]� ��������U��Vh��h�   hD ���vA  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh��h�   hD ���)A  ����t���   ��t��^��3�^����������������VW��3����$    �h��jphD ��@  ����t�@p��t	VW�Ѓ������8 tF��_��^�������U��SW��3�V��    h��jphD �@  ����t�@p��t	WS�Ѓ������8 tqh��jphD �]@  ����t�@p��t�MWQ�Ѓ�������h��jphD �+@  ����t�@p��t	WS�Ѓ�����V���������tG�]����E^��t�8��~=h��jphD ��?  ����t�@p��t	WS�Ѓ������8 u_�   []� _3�[]� ����������U��Vh��j\hD ���?  ����t3�@\��t,V��h��jxhD �g?  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh��j\hD ���)?  ����t3�@\��t,V��h��jdhD �?  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh��j\hD ����>  ����tG�@\��t@V�ЋEh��jdhD �E��E�    �E�    �>  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��j\hD ���I>  ����t\�@\��tUV��h��jdhD �'>  ����t�@d��t
�MQV�Ѓ�h��jhhD ��=  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh��j\hD ���=  ������   �@\��t~V��h��jdhD �=  ����t�@d��t
�MQV�Ѓ�h��jhhD �j=  ����t�@h��t
�URV�Ѓ�h��jhhD �A=  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh��jthD ���=  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h��j`hD ��<  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�����_�����^��]� ������U���Vh��h�   hD �u<  ����tU���   ��tK�M�UQR�M�Q�Ћu��P������h��j`hD �7<  ����t%�@`��t�U�R�Ѓ���^��]ËE�uP���k�����^��]�����U���Vh��h�   hD ����;  ����tR���   ��tH�MQ�U�R���ЋuP������h��j`hD �;  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    �'�����^��]� �������������̸   � ��������� �������������� �������������� �������������3�� �����������3�� ������������ �������������� ������������̸   � ��������3�� �����������U����E��P�X]� ������������U����E��P�X]� ������������U����E��P�X]� ������������� ������������̃��� ���������̃��� ����������3�� �����������3�� �����������3�� ����������̸   � ��������U��`��P�B<��   V�uW���Ћ}��tj VW��������u_^��]�h   ������j Q��U  �U$�E�MR�UPj QR������P�E����E�M h   ������RPWj�M��E�� �E�0� �E��� �E�`� �E�p� �E��� �E� � �E�p� �E��� �E�Э �E��� �E�� �E�@� �E��� �E��� �E�� �E�P� �EĠ� �EȰ� �E� � �q����8_^��]��̋�`L����������̋�`\����������̋�`l����������̋�`|����������̋���   �������̋�`P����������̋�``����������̋�`p����������̋���   �������̋���   �������̋�`D����������̋�`T����������̋�`d����������̋�`t����������̋���   �������̋�`H����������̋�`X����������̋�`h����������̋�`x����������̋���   ��������U��E��u�E�M�������   ]� �����������U��EHV����   �$�� �   ^]á��@�����uT�EP�k����=�2  }�����^]Ëu��t�hjmh��j���������t ���-��������tV���<����   ^]����    �   ^]ËM�UQR�b���������H^]�^]��`���-��u.�Rb���=��������t��謇��V���������    �   ^]Ã��^]ÍI  � �� �� �� ߯ ~� U��`����   �BXQ�Ѓ���u]� �`��Q|�M�RQ�MQP�҃�]� ���U��`����   �BXQ�Ѓ���u]� �`��Q|�M�R8Q�MQP�҃�]� ���U��EV��j ��`��Qj j P�B�ЉF����^]� ��̡`�Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� �`��Q�MP�EP�Q�JP�у��F�   ^]� ���̡`��H���   ��U��`��H���   V�u�R�Ѓ��    ^]����������̡`��P���   Q�Ѓ�������������U��`��P�EPQ���   �у�]� ̡`��H�������U��`��H�AV�u�R�Ѓ��    ^]��������������U��`��H�AV�u�R�Ѓ��    ^]��������������U��`��P��Vh�  Q���   �E�P�ы`����   �Q8P�ҋ�`����   ��U�R�Ѓ���^��]��������������̡`��P�BQ�Ѓ����������������U��`��P�EPQ�J\�у�]� ����U��`��P�EP�EP�EP�EP�EPQ���   �у�]� �U��`��P�EP�EP�EP�EPQ�JX�у�]� �������̡`��P�B Q��Y�U��`��P�EP�EP�EP�EPQ���   �у�]� �����U��`��P�EP�EP�EPQ�J�у�]� ������������U��`��H��   ]��������������U��`��P�R$]�����������������U��`��P��x  ]�������������̡`��P��|  ��U��`��P�EP�EP�EP�EPQ�J(�у�]� ��������U��`��P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U��`��P�EP�EP�EP�EPQ�J,�у�]� ��������U��`�V��H�QWV�ҋ��`��H�QV�ҋ`��Q�M�R4Q�MQ�MQOWHPj j V�҃�(_^]� ���������������U��`��P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U��`��P�EP�EPQ�J@�у�]� U��`��P�EPQ�JD�у�]� ���̡`��P�BLQ�Ѓ���������������̡`��P�BLQ�Ѓ���������������̡`��P�BPQ�Ѓ����������������U��`��P�EPQ�JT�у�]� ����U��`��P�EPQ�JT�у�]� ����U��`��P�EP�EPQ���   �у�]� �������������U��`��P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �`����   j P�BV�Ћ`����   �
�E�P�у� ��^��]� ������̡`��P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡`��H�������U��`��H�AV�u�R�Ѓ��    ^]��������������U��`��P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U��`��P�EPQ�J�у�]� ���̡`��P�BQ��Y�U��`��P�EP�EPQ�J�у�]� U��VW���$����M�U�x@�EPQR�������H ���_^]� �U��VW��������M�U�xD�EPQR���ޱ���H ���_^]� �V���ȱ���xH u3�^�W��趱���΍xH謱���H �_^�����U��V��蕱���xL u3�^]� W��耱���M�U�xL�EPQR���j����H ���_^]� �������������U��V���E����xP u���^]� W���/����M�U�xP�EP�EQRP�������H ���_^]� ��������U��V��������xT u���^]� W���߰���M�xT�EPQ���Ͱ���H ���_^]� U��V��走���xX u���^]� W��蟰���xX�EP��葰���H ���_^]� ����U���S�]VW���t.�M���������_����xL�E�P���Q����H ��ҍM�� ����}��tZ�`��H�A�U�R�Ћ`��Q�J�E�WP�ы`��B�P�M�Q�҃���������@@��t�`��QWP�B�Ѓ�_^[��]� ������U��V���ů���x` u
� }  ^]� W��譯���x`�EP��蟯���H ���_^]� ��U��VW��脯���xH�EP���v����H ���_^]� ���������U��SVW���S����x` u� }  �#���?����x`�E���P���,����H ��ҋ��`��H�]�QS�҃�;�A�`��H�QS�҃�;�,�������M�U�xD�EPQSR���خ���H ���_^[]� _^�����[]� ��������������U��V��襮���xP u
�����^]� W��荮���M�U�xP�EP�EQ�MR�UPQR���k����H ���_^]� ��������������U��V���E����xT u
�����^]� W���-����M�xT�EPQ�������H ���_^]� ��������������U��V��������xX tW�������xX�EP���٭���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��*  ����t.�E�;�t'�`��J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡`��H��   ��U��`��H��$  V�u�R�Ѓ��    ^]�����������U��`��UV��H��(  VR�Ѓ���^]� �����������U��`��P�EQ��,  P�у�]� �U��`��P�EQ��,  P�у����@]� �����������̡`��H��0  ��`��H��4  ��`��H��p  ��`��H��t  ��U��E��t�@�3��`��RP��8  Q�Ѓ�]� �����U��`��P�EPQ��<  �у�]� �U��`��P�EP�EP�EPQ��@  �у�]� ���������U��`��P�EP�EPQ��D  �у�]� �������������U��`��P�EPQ��H  �у�]� �U��`��P�E��L  ��VWPQ�M�Q�ҋu���`��H�QV�ҡ`��H�QVW�ҡ`��H�A�U�R�Ѓ�_��^��]� ��������������̡`��P��T  Q�Ѓ�������������U��`��P�EPQ��l  �у�]� ̡`��P��P  Q�Ѓ�������������U��`��P�EPQ��X  �у�]� ̡`��H��\  ��U��`��H��`  V�u�R�Ѓ��    ^]�����������U��`��P�EP�EP�EP�EP�EPQ��d  �у�]� �U��`��P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���2v����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���o����xP t$S���a���j j �XPj�FP���M����H ���[�    �~` t�`��H�V`�AR�Ѓ��F`    _^������������U��SV��Fx�`��Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�Tb������u#���hP�`��H��0  h  �҃��E�~P����x���j j jW�����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    �`��Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��i����F|��u�E�~x��t�    �F`_^]� �M�Fx������t�3�_^]� U��QVW�}�����&  �`��H�QhV�҃����`�u"�H��0  hPh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���$  �EF;u�|�UR�ͬ����_�   ^��]� �������������U��QVW�}����.&  �`��H�QhV�҃����`�u"�H��0  hPh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'���`��QP�Bh�Ѓ���t�M��R����#  F;u�|ʍEP������_�   ^��]� �������������hPh�   h��h�   路������t�������3��������V���(����N^��r�����������������U��VW�}�7��t��������N�r��V蝮�����    _^]á`��HL���   ��U��`��H@�AV�u�R�Ѓ��    ^]�������������̡`��HL�������U��`��H@�AV�u�R�Ѓ��    ^]�������������̡`��PL���   Q�Ѓ�������������U��`��PL�EP�EPQ���   �у�]� �������������U��`�V��HL���   V�҃���u�`��U�HL���   j RV�Ѓ�^]� �`����   �ȋBP�Ћ`����   �MP�BH��^]� �����̡`��PL��(  Q�Ѓ�������������U��`��PL�EP�EPQ��,  �у�]� ������������̡`��HL�Q�����U��`��H@�AV�u�R�Ѓ��    ^]��������������U��`��PL�E�R��VPQ�M�Q�ҋu��P���%����M��=�����^��]� ����U��`��PL�EPQ���   �у�]� �U��`��PL�EP�EPQ�J�у�]� �`��PL�BQ�Ѓ���������������̡`��PL�BQ�Ѓ���������������̡`��PL�BQ�Ѓ����������������U��`��PL�EP�EP�EPQ�J �у�]� ������������U��`��PL�EPQ��4  �у�]� �U��`��PL�EP�EP�EPQ�J$�у�]� ������������U��`��PL�EP�EP�EP�EPQ�J(�у�]� �������̡`��PL�B,Q�Ѓ���������������̡`��PL�B0Q�Ѓ����������������U��`��PL�EP�EPQ��  �у�]� ������������̡`��PL���   Q�Ѓ�������������U��`��PL�E��  ��VPQ�M�Q�ҋu��P�������M�������^��]� ̡`��PL�B4Q�Ѓ���������������̡`��PL�B8j Q�Ѓ��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL��l  ]��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL���   ]��������������U��`��PL�EPQ�J<�у�]� ���̡`��PL�BQ��Y�U��`��PL�EP�EPQ�J@�у�]� U��`��PL�Ej PQ�JD�у�]� ��U��`��PL�Ej PQ�JH�у�]� ��U��`��PL�EjPQ�JD�у�]� ��U��`��PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��t���W�M�Q�U�R���(  ���M����g�����t�`����   ��U�R�Ѓ�_^3�[��]Ë`����   �J8�E�P�ы`������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ����j�M�Q�U�R���}'  �M������`����   ��U�R�Ѓ�^��]�����������U���$�`��UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��:���j�E�P�M�Q����&  �M��1����`����   ��M�Q�҃�_^��]� ��U���$�`��UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}�����j�E�P�M�Q���y&  �M������`����   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��T���W�M�Q�U�R����%  ���M����G�����t+�u���h���`����   ��U�R�Ѓ�_��^[��]� �`����   �JL�E�P�ыu��P���%i���`����   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���4%  ���M���������t+�u����g���`����   ��U�R�Ѓ�_��^[��]� �`����   �JL�E�P�ыu��P���eh���`����   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R���t$  ���M��������_^��[t�`����   ��U�R�������]Ë`����   �J<�E�P���]��`����   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��$���W�M�Q�U�R����#  ���M���������t�`����   ��U�R�Ѓ�_^3�[��]Ë`����   �J8�E�P�ы`������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��t���W�M�Q�U�R���#  ���M����g�����t-��u�`�����   ���^�U�R�Ѓ�_��^[��]� �`����   �JP�E�P�ы�u�H��P�@�N�`��V���   �
�F�E�P�у�_��^[��]� �����̡`��PL���   Q��Y��������������U��`��PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U��`��PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R���!  ���M����������t-��u�`�����   ���^�U�R�Ѓ�_��^[��]� �`����   �JP�E�P�ы�u�H��P�@�N�`��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���   ���M���������t-��u�`�����   ���^�U�R�Ѓ�_��^[��]� �`����   �JP�E�P�ы�u�H��P�@�N�`��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��D���W�M�Q�U�R����  ���M����7�����t-��u�`�����   ���^�U�R�Ѓ�_��^[��]� �`����   �JP�E�P�ы�u�H��P�@�N�`��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��t���W�M�Q�U�R���  ���M����g�����t�`����   ��U�R�Ѓ�_^3�[��]Ë`����   �J8�E�P�ы`������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ����j�M�Q�UR���~  �M�����`����   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��O���j�U�R�E�P���  �M��F����`����   �
�E�P�у�^��]� ��������U���$�`��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}������j�E�P�M�Q���  �M�������`����   ��M�Q�҃�_^��]� ��U���$�`��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J���j�E�P�M�Q���	  �M��A����`����   ��M�Q�҃�_^��]� ��U���$�`��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}������j�E�P�M�Q���  �M�������`����   ��M�Q�҃�_^��]� ��U���$�`��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J���j�E�P�M�Q���	  �M��A����`����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E������j�U�R�E�P���  �M�������`����   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��t���W�M�Q�U�R���  ���M����g�����t-��u�`�����   ���^�U�R�Ѓ�_��^[��]� �`����   �JP�E�P�ы�u�H��P�@�N�`��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���D  ���M���藿����t�`����   ��U�R�Ѓ�_^3�[��]Ë`����   �J8�E�P�ы`������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R���  ���M���������t�`����   ��U�R�Ѓ�_^3�[��]Ë`����   �J8�E�P�ы`������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ���̡`��PL���  ��U���$�`��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}������j�E�P�M�Q���  �M������`����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�����j�U�R�E�P���N  �M�膽���`����   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�����j�U�R�E�P����  �M������`����   �
�E�P�у�^��]� ��������U��`��H���   ]��������������U��`��H���   ]�������������̡`��H���   ��`��H���   ��U��`��H���   V�u�R�Ѓ��    ^]�����������U��`��H���   ]��������������U��`��HL�QV�ҋ���u^]á`��H�U�Ej R�UP��h  RV�Ѓ���u�`��Q@�BV�Ѓ�3���^]��������U��`��H�U�E��h  j R�U�� P�ERP�у�]����U��`��H���   ]��������������U��`��H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡`��PL�BLQ�Ѓ���������������̡`��PL�BPQ�Ѓ����������������U��`��PL�EP�EPQ�JT�у�]� U��`��PL�EPQ��  �у�]� �U��`��PL�EPQ���   �у�]� ̡`��PL�BXQ�Ѓ����������������U��`��PL�EP�EP�EPQ�J\�у�]� ������������U���4�`�SV��HL�QW�ҋ�3ۉ}�;��x  �M������`��E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ`����   �BSSW���Ѕ���   �`��QL�BW�Ћ���;���   ��    �`����   �B(���ЍM�Qh�   ���u��A��������   �M�;���   �`����   ���   S��;�tm�`����   �ȋB<V�Ћ`����   ���   �E�P�у�;�t�`��B@�HV�у���;��\����}��M���U���M�������_^[��]� �}��`��B@�HW�ы`����   ���   �M�Q�҃��M��yU���M��ѵ��_^3�[��]� �����̡`��PL�B`Q�Ѓ���������������̡`��PL�BdQ�Ѓ����������������U��`��PL�EPQ�Jh�у�]� ���̡`��PL��D  Q�Ѓ������������̡`��PL�BlQ�Ѓ����������������U��`��PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh`� h@� h � h� R�Q�U R�UR�UR�U���A�$�5`��vLRP���   Q�Ѓ�4^]�  ������̡`��PL���   Q�Ѓ�������������U��`��PL�EP�EP�EPQ��   �у�]� ���������U��`��PL��H  ]�������������̡`��PL��L  ��U��`��PL��P  ]��������������U��`��PL��T  ]��������������U��`��PL��p  ]��������������U��`��PL��t  ]��������������U��`��PL�EP�EP�EP�EP�EPQ���   �у�]� �U��`��PL�EP�EP�EPQ���   �у�]� ���������U��`��PL�EP�EP�EP�EPQ��   �у�]� �����U��`��HL���   ]��������������U��`��HL���   ]��������������U��`��HL���   ]�������������̡`��HL��  ��`��HL��@  ��U��`��PL���  ]��������������U��`��PL���  ]��������������U��`��PL���  ]��������������U��� �`�V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�`��QLjP���   ���ЋM��U�Rh=���M�}��S<�����`����   ���   �U�R�Ѓ��M��u���P����_^��]Ë`����   ���   �E�P�у��M��u��P��_�   ^��]����U��� �`�V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�`��QLjP���   ���ЋM��U�Rh<���M�}��;�����`����   ���   �U�R�Ѓ��M��u���O����_^��]Ë`����   ���   �E�P�у��M��u���O��_�   ^��]����U��E�M�UP��P�EjP��=����]��������������̸   �����������U��V�u��t���u6�EjP��=������u3�^]Ë���>����t���t��U3�;P��I#�^]�������h��Ph�f �������������������U��h��jh�f �|�������t
�@��t]�����]�������U��Vh��jh�f �K���������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�P���E�NP�у�4�M���DP����^]ÍM�7P�����^]��U��h��jh�f ���������t
�@��t]��3�]��������U��h��jh�f ��������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á`��H�F��  h�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�c���3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�A�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W���m���3����_�F�F^��������������U���SV�uW���^S�}��6���3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY�`��H���  h�j8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E���K  ��]� �����U����Q�Ej�E��A�MRPQ�M��E���g  ��]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q����t!�A��t�B�A�Q�P�A    �A    �̋�� ��@��HV3��q�q�P�r�r���p�p�p�P�H^������V���������F3��F�;�t�N;�t�H�F�N�H�V�V�F�F�;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3���;�t�F;�t�A�F�N�H�V�V�Et	V�&�������^]� ������������U��V��W�~W��躀��3����E��F�Ft	V������_��^]� ������U��V��������Et	V蹃������^]� ��������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�`����   P�B@��]� �E��t�`����   P�BD��]� �`����   R�PD��]� �����U��`��P@�Rd]�����������������U��`��P@�Rh]�����������������U��`��P@�Rl]�����������������U��`��P@�Rp]�����������������U��`����   ���   ]�����������U��`����   ���   ]����������̡`��P@�Bt����̡`��P@�Bx�����U��`��P@�R|]����������������̡`��P@���   ��`����   �Bt��U��`��P@���   ]�������������̡`��P@���   ��U��`��P@���   ]��������������U��`��P@���   ]��������������U��`��P@���   ]��������������U��`��P@���   ]��������������U��`��P@���   ]��������������U��`��P@���   ]��������������U��`�V��H@�QV�ҋM����t��#����`��Q@P�BV�Ѓ�^]� �̡`��PH���   Q�Ѓ�������������U��`��P@�EPQ�JL�у�]� ���̡`��P@�BHQ�Ѓ����������������U��`��P@�EP�EP�EPQ�J�у�]� ������������U��`��P@�EPQ�J�у�]� ����U��`��P@�EP�EPQ�J�у�]� U��`��P@�EPQ�J �у�]� ����U��`����   �R]��������������U��`����   �R]��������������U��`����   �R ]��������������U��`����   ���   ]�����������U��`����   ��D  ]�����������U��`��E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U��`����   ���   ]����������̡`����   �B$��`��H@�Q0�����U��`��H@�A4j�URj �Ѓ�]����U��`��H@�A4j�URh   @�Ѓ�]�U��`��H@�U�E�I4RPj �у�]�̡`��H|�������U��V�u���t�`��Q|P�B�Ѓ��    ^]��������̡`��H|�Q �����U��V�u���t�`��Q|P�B(�Ѓ��    ^]��������̡`��H@�Q0�����U��V�u���t�`��Q@P�B�Ѓ��    ^]���������U��`��H@���   ]��������������U��V�u���t�`��Q@P�B�Ѓ��    ^]��������̡`��PH���   Q�Ѓ�������������U��`��PH�EPQ��d  �у�]� �U��`��H �IH]�����������������U��}qF uHV�u��t?�`����   �BDW�}W���Ћ`��Q@�B,W�Ћ`��Q�M�Rp��VQ����_^]����������̡`��P@�BT�����U��`��P@�RX]�����������������U��`��P@�R\]����������������̡`��P@�B`�����U��`��H��T  ]��������������U��`��H@�U�A,SVWR�Ћ`��Q@�J,���EP�ы`��Z��h��hE  �΋�薟��Ph��hE  ��脟��P��T  �Ѓ�_^[]����U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� ø*����������� �g�$��(���,���0���4�rË�U�������4  �} ���t�  ��]�;p�u���
  ��Q��  YË�U��V��������EtV�qt��Y��^]� ��U��EVW��u|P�!0  Y��u3��  �9#  ��u�70  ���/  �����m.  ����(  ��}�  ���-  ��| �+  ��|j �F&  Y��u����   �*  ��3�;�u19=��~����9=T�u��'  9}u{�|*  �P  �/  �j��uY�  h  j�Y$  ��YY;��6���V�5@��5��f  Y�Ѕ�tWV�D  YY� �N���V�  Y�������uW��!  Y3�@_^]� jh ��1  ����]3�@�E��u9����   �e� ;�t��u.���tWVS�ЉE�}� ��   WVS�r����E����   WVS�����E��u$��u WPS����Wj S�B������tWj S�Ѕ�t��u&WVS�"�����u!E�}� t���tWVS�ЉE��E������E���E��	PQ�$0  YYËe��E�����3��x0  Ë�U��}u�
2  �u�M�U�����Y]� ��U��QSVW�5����  �5�����}���  ��YY;���   ��+ߍC��rwW�K2  ���CY;�sH�   ;�s���;�rP�u���"  YY��u�G;�r@P�u��"  YY��t1��P�4��  Y����u��  ���V��  Y����EY�3�_^[�Ë�Vjj �"  ��V��  ����������ujX^Ã& 3�^�jh@��/  �#  �e� �u�����Y�E��E������	   �E��4/  ���"  Ë�U���u���������YH]�������������̋T$�L$��ti3��D$��u��   r�=�� t�2  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh`��>.  �e� �u;5��w"j�j4  Y�e� V�q<  Y�E��E������	   �E��J.  �j�e3  YË�U��V�u�����   SW�=�=l� u�@  j�?  h�   �!  YY�����u��t���3�@P���uV�S���Y��u��uF�����Vj �5l��׋؅�u.j^9��t�u� A  Y��t�u�{����@  �0�@  �0_��[�V��@  Y�@  �    3�^]�jh���%-  �u��tu�=��uCj�P3  Y�e� V�x3  Y�E��t	VP�3  YY�E������   �}� u7�u�
j�<2  Y�Vj �5l����u�@  ���P��?  �Y��,  ���������������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�i@  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�@  ���$�2D  �   ��ÍT$��C  R��<$tPf�<$t�-8&������z�=�� �D  �   ����	D  �-:&��������z��������oC  ���� u�|$ u����-��   �=�� ��C  �   ����D  Z�������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��D  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�uD  ���$�C  �   ��ÍT$�B  R��<$tPf�<$t�-8&������z�=�� ��B  �   �����B  �-:&��������z��������?B  ���� u�|$ u����-��   �=�� ��B  �   ����C  Z�������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�IE  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u��D  ���$��A  �   ��ÍT$�}A  R��<$t6f�<$t�-8&����=�� ��A  �   ����A  �)A  �&��� u�|$ u����-���   �t���뻸   �=�� �fA  �   ����_B  Z������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�G  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u��F  ���$�@  �   ��ÍT$�]@  R��<$tL�D$f�<$t�-8&�  �t^�   �uA������=�� �|@  �б�   �y@  �   �u�ԩ�� u�|$ u%   �t����-��   �"��?  ���� uŃ|$ u����-*��   �=�� �@  �б�   �	A  ZÃ��$��?  �   ��ÍT$�?  R��<$�D$tQf�<$t�@?  �   �u���=�� ��?  �   ���?  �  �u,��� u%�|$ u���?  �"��� u�|$ u�%   �t����-��   �=�� �V?  �   ���O@  Z������̃=�� �JL  ���\$�D$%�  =�  u�<$f�$f��f���d$�L  � �~D$f(0f(�f(�fs�4f~�fT`f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$��H  ���D$��~D$f��f(�f��=�  |!=2  �fT �\�f�L$�D$����f�PfVPfT@f�\$�D$���������������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��K  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�K  ���$�r=  �   ��ÍT$�=  R��<$tmf�<$t��<  =  �?s+��������������=�� �@=  �   ���==  w:�D$��%�� D$u)��   ����-��t�����<  ���� u�|$ u����-��   �=�� ��<  �   ����=  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�	P  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�O  ���$�"<  �   ��ÍT$��;  R��<$tmf�<$t�;  =  �?s-����������������=�� ��;  �   � ���;  w8�D$��%�� D$u'��   ���t��������B;  ���� u�|$ u����-��   �=�� ��;  �   � ��<  Z����������̺���aU  �����T  �����������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�Ë�U��EV���F ��uc�  �F�Hl��Hh�N�;�t���Hpu�Ta  ��F;�t�F���Hpu��Y  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P�Td  ��e�F�P�c  ��Yu��P�7d  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�sc  �M��E��M��H��EP�d  �E�M����Ë�U��j �u�u�u������]Ë�V����tV��g  @PV�V�wd  ��^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+�l3  j_VVVVV�8��`  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�(3  j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]hpSV�ag  ��3ۅ�tSSSSS��^  ���N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�8�t�90uj�APQ��b  ���}� t�E��`p�3�_^[�Ë�U���,�p�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�h  3ۃ�;�u��1  SSSSS�0�N_  �����o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�f  ��;�t���u�E�SP�u��V�u��������M�_^3�[�V����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �C���9}}�}�u;�u+��0  j^WWWWW�0�a^  ���}� t�E�`p����  9}vЋE��� 9Ew	�0  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�4R  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� �Lg  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� ��f  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���WF�f  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP�_e  0�F�U�����;�u��|��drj jdRP�9e  0��U�F����;�u��|��
rj j
RP�e  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�������u-�-  j^�03�PPPPP��Z  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�������}� t�E��`p�3�_^[�Ë�U���,�p�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�,c  3ۃ�;�u�,  SSSSS�0��Y  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P�Za  ��;�t���u�E�SV�u���`������M�_^3�[�����Ë�U���0�p�3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�qb  3ۃ�;�u��+  SSSSS�8�9Y  �����   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW�`  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�����Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3�����6�x  ��Y���(r�_^Ë�Vh   h   3�V�eb  ����tVVVVV�pV  ��^Ë�U������]��x�]��E��u��M��m��]����]�����z3�@��3���h����th�P���tj ���������U��� S3�9]u �)  SSSSS�    �W  ������   �MV�u;�t!;�u�o)  SSSSS�    ��V  ������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u���c  ����;�t�M�x�E����E�PS�a  YY��_^[�Ë�U���uj �u�u�u�5�����]Ë�U���(  �������������5���=��f��f���f���f���f�%��f�-���� ��E ����E����E���������@�  ���������	 ����   �p��������t��������,�8�j�Yn  Yj �(h��$�=8� uj�5n  Yh	 �� P���jh���r  j�  Y�e� �u�N��t/�����E��t9u,�H�JP�
���Y�v����Y�f �E������
   �a  Ë���j�x  Y����������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U��V�5D��54�օ�t!�@����tP�5D����Ѕ�t���  �'��V�0��uV�  Y��th�P���t�u�ЉE�E^]�j ����YË�U��V�5D��54�օ�t!�@����tP�5D����Ѕ�t���  �'��V�0��uV�   Y��th�P���t�u�ЉE�E^]��8� ��V�5D��4����u�5��e���Y��V�5D��<��^á@����tP�5 ��;���Y�Ѓ@���D����tP�@�D���&  jh���	  ��V�0��uV�a  Y�E�u�F\H3�G�~��t$h�P��Ӊ��  h��u��Ӊ��  �~pƆ�   CƆK  C�Fh�j��  Y�e� �vh�D�E������>   j�  Y�}��E�Fl��u���Fl�vl�O  Y�E������   �  �3�G�uj�  Y�j�  YË�VW��5@��������Ћ���uNh  j��  ��YY��t:V�5@��5������Y�Ѕ�tj V�����YY� �N���	V����Y3�W�H_��^Ë�V��������uj�>  Y��^�jh��  �u����   �F$��tP�F���Y�F,��tP�8���Y�F4��tP�*���Y�F<��tP����Y�F@��tP����Y�FD��tP� ���Y�FH��tP�����Y�F\=HtP�����Yj�L  Y�e� �~h��tW�L��u���tW����Y�E������W   j�  Y�E�   �~l��t#W�N  Y;=�t���t�? uW�L  Y�E������   V�\���Y��  � �uj��  YËuj��  YË�U��=@��tK�} u'V�5D��54�օ�t�5@��5D����ЉE^j �5@��5�����Y���u�x����D����t	j P�<]Ë�VW��V�0��uV�R  Y�����^  �5hW��hW����h�W����h�W���փ=� �5<� �t�=� t�=� t��u$�4���@����5�� ��8�D������   �5�P�օ���   �_  �5������5��������5��������5 ����u������ ��  ��teh� �5������Y�У@����tHh  j�   ��YY��t4V�5@��5�����Y�Ѕ�tj V�y���YY� �N��3�@��$���3�_^Ë�U��VW3��u�e�����Y��u'9$�vV�P���  ;$�v��������uʋ�_^]Ë�U��VW3�j �u�u�h  ������u'9$�vV�P���  ;$�v��������uË�_^]Ë�U��VW3��u�u��h  ��YY��u,9Et'9$�vV�P���  ;$�v��������u���_^]Ë�U��W��  W�P�u�0���  ��`�  w��t�_]Ë�U���<  �u�  �5H��D���h�   �Ѓ�]Ë�U��h0�0��th P���t�u��]Ë�U���u�����Y�u�T�j�1  Y�j�N  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=  th �Wj  Y��t
�u� Y�p���h@h(����YY��uBh/�p�����$$�c����=�� Yth����i  Y��tj jj ���3�]�jh��  j�M  Y�e� 3�C9X���   �T��E�P��} ��   �5�������Y���}؅�tx�5������Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5���~������5���q�����9}�u9E�t�}�}؉E����u܋}��hP�D�_���YhX�T�O���Y�E������   �} u(�X�j�{  Y�u�����3�C�} tj�b  Y��8
  Ë�U��j j�u�������]�jj j ������Ë�V������V�e  V�k  V�RI  V��>  V�k  V�ri  V�x���V�Ui  hb'������$�H�^�jTh0��s	  3��}��E�P�d�E�����j@j ^V�&���YY;��  ����5����   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�����   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M��������� ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=��|���=���e� ��~m�E����tV���tQ��tK�uQ�`��t<�u���������4����E� ���Fh�  �FP�
j  YY����   �F�E�C�E�9}�|�3ۋ���5������t���t�N��r�F���uj�X�
��H������P�\�����tC��t?W�`��t4�>%�   ��u�N@�	��u�Nh�  �FP�ti  YY��t7�F�
�N@�����C���g����5���X3��3�@Ëe��E���������q  Ë�VW����>��t1��   �� t
�GP�h���@   ;�r��6�����& Y������|�_^Ã=�� u�-C  V�5��W3���u����   <=tGV�:N  Y�t���u�jGW�n�����YY�=8���tˋ5��S�BV�	N  ��C�>=Yt1jS�@���YY���tNVSP�sN  ����t3�PPPPP��E  �����> u��5��� ����%�� �' ���   3�Y[_^��58�������%8� ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�[h  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�vg  Y��t��M�E�F��M��E���Sg  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9��u�@  h  �`�VS�d��l����5H�;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�q�����Y;�t)�U��E�P�WV�}�������E���H�,��50�3�����_^[�Ë�U��h���SV�5�W3�3�;�u.�֋�;�t�h�   �#���xu
jX�h���h�����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5|SSS+�S��@PWSS�E��։E�;�t/P����Y�E�;�t!SS�u�P�u�WSS�օ�u�u�����Y�]��]�W�x���\��t;�u��t��;��r���8t
@8u�@8u�+�@P�E��0�����Y;�uV�p�E����u�VW�`e  ��V�p��_^[�Ë�V����W��;�s���t�Ѓ�;�r�_^Ë�V����W��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P���l���u]�3�@���]Ã=��uWS3�9��W�=~3V�5����h �  j �v����6j �5l��׃�C;��|�^�5��j �5l���_[�5l����%l� Ë�U��QQV�H��������F  �V\���W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ����=�����;�}$k��~\�d9 �=�����B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]����h�1d�5    �D$�l$�l$+�SVW�p�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���̋�U���S�]V�s35p�W��E� �E�   �{���t�N�38������N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���Y  �E���|@G�E��؃��u΀}� t$����t�N�38�K����N�V�3:�;����E�_^[��]��E�    �ɋM�9csm�u)�=�� t h���s]  ����t�UjR������M�WY  �E9Xthp�W�Ӌ��ZY  �E�M��H����t�N�38�����N�V�3:�����E��H����X  �����9S�R���hp�W���Y  ������U����p��e� �e� SW�N�@��  ��;�t��t	�Уt��`V�E�P���u�3u���3�� 3���3��E�P���E�3E�3�;�u�O�@����u������5p��։5t�^_[��jhP��v���3��]3�;���;�u��  �    WWWWW�)>  ������S�=��u8j�{  Y�}�S�  Y�E�;�t�s���	�u���u��E������%   9}�uSW�5l��������6����3��]�u�j�I  Y�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jhp�������e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E������Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[���������3�Ë�VW3��p��<���u�����8h�  �0���]  YY��tF��$|�3�@_^Ã$��� 3����S�hV���W�>��t�~tW��W�����& Y����ȳ|ܾ��_���t	�~uP�Ӄ���ȳ|�^[Ë�U��E�4Ũ���]�jh���u���3�G�}�3�9l�u�D  j�  h�   �A���YY�u�4���9t���nj�����Y��;�u�  �    3��Qj
�Y   Y�]�9u,h�  W�\  YY��uW�����Y�Q  �    �]���>�W����Y�E������	   �E������j
�(���YË�U��EV�4Ũ��> uP�"���Y��uj�5���Y�6��^]Ë�U�������k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �������   ����5�h @  ��H� �  SQ�֋������   ���	P����@�������    ����@�HC����H�yC u	�`�����x�ueSj �p�֡���pj �5l��������k����+ȍL�Q�HQP�:  �E�����;��v�m�������E����=��[_^�á��V�5��W3�;�u4��k�P�5��W�5l���;�u3��x����5�����k�5��h�A  j�5l���F;�t�jh    h   W���F;�u�vW�5l��뛃N��>�~����F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W����u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U�������Mk���������M���SI�� VW}�����M���������3���U��������S�;#U�#��u
���];�r�;�u�����S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1����	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t����C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;��u�M�;��u�%�� �M���B_^[�Ë�U��QQS�]VW3�3��}�;�ȳt	G�}���r���w  j�dW  Y���4  j�SW  Y��u�=���  ���   �A  hh�  S���W�c6  ����tVVVVV��-  ��h  ���Vj ��� �l��u&hPh�  V�!6  ����t3�PPPPP�-  ��V�z5  @Y��<v8V�m5  ��;�j���hL+�QP��U  ����t3�VVVVV�d-  ���3�hHSW�KU  ����tVVVVV�@-  ���E��4�̳SW�&U  ����tVVVVV�-  ��h  h W�S  ���2j��\��;�t$���tj �E�P�4�̳�6�4  YP�6S��_^[��j��U  Y��tj��U  Y��u�=��uh�   �)���h�   ����YYË�U��E3�;̀�tA��-r�H��wjX]Ë̈́�]�D���jY;��#���]��n�����u��Ã���[�����u��Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E���]Ë�U���5���8���Y��t�u��Y��t3�@]�3�]Ã%�� �l������3�����������U�������$�~$�   ��fD$f��f%�f-00f=��B  f�%�Y�f�%�-��X�f�%�\�f(�%�Y�fɁ� v ����?f(-�%�����fY��\��Y�%�\�fxf����\�fY�f\�f(5�%�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�%�Y fX5�%fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y&fD$�D$���f &�Y��\��Y&fD$�D$����8�����������̀zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp��������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-���p��� ƅp���
��
�t�����������������������������ËT$��   ��f�T$�l$é   t�   ��0&�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ��   Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�{   Z��]   Z��,$Z��\&�����������L&�����   s��l&��T&�����������D&�����   v��d&�����U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�O  ���E�f�}t�m���������������U�������$�~$�   ��fD$f��f%�f-00f=��B  f�.�Y�f�.�-��X�f�.�\�f(�.�Y�fɁ�v ����?f(-�.��&���fY��\��Y�.�\�fxf����\�fY�f\�f(5�.�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�.�Y fX5�.fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f/�\�fL$�D$���������I ����U�������$�~<$�   ���~|$f�f(�fT@/f/h0��  �U  f/X0snf/`0��  f(�fY�f(�fY�f(-0fY�fX- 0fY�fX-�/fY�fX-�/�Y�f(�f���X��Y��\�f�|$�D$�f/P0��   f(�fY�f(�fY�f(-�/fY�fX-�/fY�fX-�/fY�fX-�/fY�fX-�/fY�fX-�/fY�fX-p/fY�fX-`/�Y�f(�f���X��Y��\�f�|$�D$��~�fW�f/H0sO�~@0�~- 0�~��X�fs�,f��f~؍@�~,�s�~��\��Y��X80�^�f���   �~��~00�^�f��~��r�~$� sf(�fY�f(�fY�f(-0fY�fX- 0fY�fX-�/fY�fX-�/�Y�f(�f���X��Y��\��\��\�fV�f�D$�D$�f/(0u�D$�f/p0s�x0�x0���$�$���D$��x0�x0�D$��~��~0/fT�f.�z�D$���x0��P/ú�  ���T$�ԃ��T$�T$�$�  ���D$Ð����U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(�0f(�0f(%�0f(5�0fT�fV�fX�f�� %�  f(�`1f(�p5fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(01f(�f(@1fY�fY�fX�f(P1�Y�f(-�0fY�f(��0fT�fX�fX�fY��Y�fX�f(�f�fY˃�f(�f��X��X��X�fD$�D$���fD$f(�0��� f�� �� wH���t^���  wlfD$f(�0f(�0fT�fV���� f�� �� t�1ú�  �Of�0�^�f1�   �4f 1�Y�������/��������  ���  s:fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$�@  �D$���fT$fD$f~�fs� f~с��� ��� t���  릍d$ ƅp����
�uK�����ƅp����2������;  ������a���t��=��t����S  ��@u��
�t��������F  �t2��t�������������^��������- �ƅp����������ݽ`������a���Au����ƅp������-*��
�uS��������
�u�����n�����   ����
�u���u
�t���ƅp����- ���u�
�t��������-����������X��ݽ`������a���u���- �
�t���ƅp�������������- �ƅp����
�u����- �������->��ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���R������ٛ���t�   ø    ���   ��V��t��V���$���$��v�6H  ���f���t^��t�����Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9��t�5������Y����M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�<:��M��]�Q��]���]���Y����  ������ "   �  �E�8:��M��]�Q��E�   �]���]���Y�j  �E�   �E�8:��E�0:��]���]���"  �M��E�0:�r����E�,:�׉M��E�,:�Z����E�<:놃�tNIt?It0It ��t����   �E�$:��E�:��E�<:����E�<:�x����E�   ��������   �E�   �E�:��������������   �$�sV�E�,:��E�0:��E�8:��E�:��E�:��E��9�y����E��9�m����E��9��E��9��E��9��M����]���]�M��]�Q�E�   ��Y��u�P���� !   �E��_^[���U�U�U�U�UV�UV|UsUV(V1V��U��QQSV���  V�5|��\  �EYY�M�ظ�  #�QQ�$f;�uU�M[  YY��~-��~��u#�ESQQ�$j��Y  ���rVS�[\  �EYY�d�ES�����\$�E�$jj�?�Z  �]��EY�]�Y����DzVS�\  �E�YY�"�� u��E�S���\$�E�$jj�Y  ��^[������U�������$�~$�   ��fD$f%�Qf�QfW�f�Q��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fUPIfV�f($�P:���X��\��Y��Y��Y����X��^�f=�Qf-�Q�\�fs�?��fs�?�Y�fp�Df5�Q�Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT=�Qfs���f%�Q���\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<�PI�Y�f(PQ�Y��Y��\��X��\��X�f-�Q�\��X�f�Q�^�f�Qf\�P:���Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5�Qf�f(�Qf(%�QfY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=pQfp�DfTpQ��f%�Q���\��Y��X��Y��\����Y��Y��\��\��X��\�f(�Qfp���\��X�fp���X��Y��X�fp���^�f(�Qf(-�Qf(�QfY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(PQ�Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$����fD$����fD$�D$���f�QfPQfXQ�X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$���U�������$�~$�   ��fD$f%�if jfW�f�i��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU0afV�f($�0R���X��\��Y��Y��Y����X��^�f�if-�i�\�fs�?��fs�?�Y�fp�Df5�i�Y��Y���fW��Y�f\%0i�Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<�0a�Y��Y��Y��\�fT@i�X��\��X�f-�i�\��X�f�i�^�f�ifX�0R���Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(5�if�f(�if(%�ifY�f(-0i��fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT=�if%jf(�i�Y�f(�i�\�f(�ifp�D�Q�fY�fp�Df��fY�fX�fpifY�����Y�fX�fp�D�Y�fT@ifY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�4���fD$����fD$�D$���f������fn�fp� fPifXifT�fT��X�fD$�D$���f0if8i�X�fD$�D$���fW��Xƺ�  �J����������������7   ���"�.   ��������2��ƅp��������������
�t����
�t�����������������������ݽ`������a���u2����X��������-�����
�t����
�t�������
�t������������؊�� ������������������U���0���S�ٽ\�����=p� t�W�����8����   [����ݕz������U���U���0���S�ٽ\����=p� t������8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq��������   [�À�8�����=�� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �Xj�����������Hj����s4�hj�,ǅr���   �Pj�����������@j����v�`jVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�^5  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�������������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Ë�U���(  �p�3ŉE��жVtj
�����Y��+  ��tj��+  Y�ж��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�1�������������(�����0���j ǅ����  @��������,����(��(���P�$j����̋�U��E���]�����������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�]���3��ȋ��~�~�~����~��������F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �p�3ŉE�SW������P�v���   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R蚚����C�C��u�j �v�������vPW������Pjj ��Q  3�S�v������WPW������PW�vS��O  ��DS�v������WPW������Ph   �vS�O  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[覕����jh���5����{��������Gpt�l t�wh��uj 讻��Y���M����j�B���Y�e� �wh�u�;5�t6��tV�L��u���tV蟚��Y���Gh�5��u�V�D�E������   뎋u�j����YË�U���S3�S�M�� ���������u���   ��8]�tE�M��ap��<���u���   ���ۃ��u�E��@���   ��8]�t�E��`p���[�Ë�U��� �p�3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9����   �E��0=�   r����  �p  ����  �d  ��P�����R  �E�PW�����3  h  �CVP躗��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�s����M��k�0�u��� ��u��*�F��t(�>����E����D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C���Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95���X�������M�_^3�[衒����jhК�0����M���r������}�������_h�u�u����E;C�W  h   苷��Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�L��u�Fh=�tP�{���Y�^hS�=D���Fp��   ����   j�����Y�e� �C���C���C��3��E��}f�LCf�E��@��3��E�=  }�L�� �@��3��E�=   }��  ���@���5��L��u��=�tP���Y��S���E������   �0j�<���Y��%���u ���tS茖��Y�����    ��e� �E������Ã=�� uj��V���Y���   3�Ë�U��SV�u���   3�W;�to=p�th���   ;�t^9uZ���   ;�t9uP�������   � N  YY���   ;�t9uP�������   �M  YY���   �ڕ�����   �ϕ��YY���   ;�tD9u@���   -�   P讕�����   ��   +�P蛕�����   +�P荕�����   肕�������   �=��t9��   uP�K  �7�[���YY�~P�E   ���t�;�t9uP�6���Y9_�t�G;�t9uP����Y���Mu�V����Y_^[]Ë�U��SV�5DW�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5LW�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu���tV�Y���Y��^�3��jh��������������Fpt"�~l t������pl��uj �=���Y��������j�����Y�e� �Fl�=��i����E��E������   ��j�����Y�u�Ë�U��E�4�]Ë�U���(  �p�3ŉE������� SjL������j P�_�����������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������,j ���(��(���P�$��u��uj��  Yh �� P��M�3�[荌���Ë�U���54�����Y��t]��j�  Y]������U����u�M�膜���E����   ~�E�Pj�u��J  ������   �M�H���}� t�M��ap��Ë�U��=� u�E�ؼ�A��]�j �u����YY]Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS�VJ  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�J  YY��t�Ej�E��]��E� Y��+���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�hD  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=� u�E�H���w�� ]�j �u�����YY]Ë�U���(�p�3ŉE�SV�uW�u�}�M�賚���E�P3�SSSSW�E�P�E�P�T  �E�E�VP�J  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������Ë�U���(�p�3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P��S  �E�E�VP�N  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�W�������������������U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�Z  ��   u������r*��$��v��Ǻ   ��r����$��u�$��v��$�xv�v4vXv#ъ��F�G�F���G������r���$��v�I #ъ��F���G������r���$��v�#ъ���������r���$��v�I �v�v�v�v�v�v�v�v�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��v���v�vww�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��x�����$�0x�I �Ǻ   ��r��+��$��w�$��x��w�w�w�F#шG��������r�����$��x�I �F#шG�F���G������r�����$��x��F#шG�F�G�F���G�������V�������$��x�I 4x<xDxLxTx\xdxwx�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��x���x�x�x�x�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��MS3�VW;�t�};�w�+���j^�0SSSSS���������0�u;�u��ڋъ�BF:�tOu�;�u������j"Y�����3�_^[]Ë�U��MSV�u3�W�y;�u�����j^�0SSSSS�.��������   9]v݋U;ӈ~���3�@9Ew����j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�a���@PWV�������3�_^[]Ë�U��Q�M�ASVW������  #�% �  �߉E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��E��<  �U����������U��E�����P������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0�p�3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��U  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�A������M�_�s^��3�[�߂����������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j����YË�U��E�M%����#�V������t1W�}3�;�tVV�^  YY�����j_VVVVV�8� �������_��uP�u��t	�^^  ���U^  YY3�^]Ë�U��QV�uV�\m  �E�FY��u�?���� 	   �N ����/  �@t�$���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�9k  �� ;�t�-k  ��@;�u�u�j  Y��uV�fj  Y�F  W��   �F�>�H��N+�I;��N~WP�u�Zi  ���E��M�� �F����y�M���t���t���������������P��@ tjSSQ��`  #����t%�F�M��3�GW�EP�u��h  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�m����8*u�ϰ?�d����} �^[]Ë�U���x  �p�3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������&�����u5������    3�PPPPP�L����������� t
�������`p������
  �F@u^V�j  Y�P����t���t�ȃ��������������A$u����t���t�ȃ������������@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw�����j��3��3�3����kj��Y������;���	  �$�֊��������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������!;  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P��g  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  � �������P����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������`e  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V讝��������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5(�觗��Y�Ћ���������   t 9�����u������PS�54��x���Y��YY������gu;�u������PS�50��S���Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�9d  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u� ��������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�wb  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t�������y�������� Y���������������t������������������������� t
�������`p��������M�_^3�[��s���Ð���p���ǁ�;��%�� ���SVW�T$�D$�L$URPQQh��d�5    �p�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�.c  �   �C�@c  �d�    ��_^[ËL$�A   �   t3�D$�H3��s��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�b  3�3�3�3�3���U��SVWj j h7�Q�t  _^[]�U�l$RQ�t$������]� jh�������M3�;�v.j�X3���;E�@u�7����    WWWWW������3���   �M��u;�u3�F3ۉ]���wi�=��uK������u�E;��w7j�ª��Y�}��u�Ȳ��Y�E��E������_   �]�;�t�uWS�u����;�uaVj�5l����;�uL9=��t3V����Y���r����E;��P����    �E���3��uj�f���Y�;�u�E;�t�    ���)����jh0��ף���]��u�u��u��Y��  �u��uS�v��Y�  �=����  3��}�����  j�ϩ��Y�}�S�����Y�E�;���   ;5��wIVSP�ڮ������t�]��5V話��Y�E�;�t'�C�H;�r��PS�u��  S訩���E�SP�Ω����9}�uH;�u3�F�u������uVW�5l���E�;�t �C�H;�r��PS�u���  S�u�聩�����E������.   �}� u1��uF������uVSj �5l�������u�]j� ���YË}����   9=��t,V�4���Y��������ε��9}�ul���P�y���Y��_����   詵��9}�th�    �q��uFVSj �5l�������uV9��t4V�˵��Y��t���v�V軵��Y�]����    3��6�����J����|�����u�<������P�����Y�������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�hP�h�1d�    P��SVW�p�1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jhp��k���豏���@x��t�e� ���3�@Ëe��E���������脠���hݐ踌��Y�x�Ë�U��E�|����������]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5���̌��Y�j h��迟��3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�e������}؅�u����a  �|��|��`�w\���]���������Z�Ã�t<��t+Ht讲���    3�PPPPP������뮾�������������
�������E�   P�����E�Y3��}���   9E�uj�����9E�tP�$���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.����M܋������9M�}�M�k��W\�D�E����p�����E������   ��u�wdS�U�Y��]�}؃}� tj 貣��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��a���Ë�U��E���]Ë�U��E���]�jh�������e� �u�u���E��/�E� � �E�3�=  �����Ëe�}�  �uj�H�e� �E������E�����Ë�U����u�M��!{���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]���������������U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]��;  ��   u������r*��$�����Ǻ   ��r����$����$�����$�8��Ȕ���#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I ������x�p�h�`�X��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������ȕܕ�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�@������$���I �Ǻ   ��r��+��$�D��$�@��T�x����F#шG��������r�����$�@��I �F#шG�F���G������r�����$�@���F#шG�F�G�F���G�������V�������$�@��I ��������$�7��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�@���P�X�h�|��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U���SVW襆���e� �=�� ����   h�r�������*  �5h�rW�օ��  P�����$�rW�����P�څ���$�rW�����P�Ņ���$�rW�����P谅��Y�����th�rW��P蘅��Y������;�tO9��tGP������5��������YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9���;�t0P覅��Y��t%�ЉE���t���;�tP艅��Y��t�u��ЉE��5���q���Y��t�u�u�u�u����3�_^[�Ë�U��ES3�VW;�t�};�w蘫��j^�0SSSSS���������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��Q���j"Y����3�_^[]Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w����j^�0SSSSS�y���������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x����蕪��j"Y���낋�U��MV3�;�|��~��u����(��������Z���VVVVV�    ����������^]Ë�S��QQ�����U�k�l$���   �p�3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|�����  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�b  ��h��  ��x�����  �>YYt�=p� uV�Z  Y��u�6�2  Y�M�_3�^�c����]��[Ë�U��QQ�EQQ�$��R  YY��uH�EQQ�$�  �]YY����Dz/�EQ��Q�]��E��$��  �]�YY����DzjX��3�@��3��Ë�U����V�U3�3����E��Au��  ��  ��9Eu=9Uu��������z�������`���   ��������A�Eu����   ����   9MuB9Uu=��������z	�����   ���������Ez�`��   �h�3��F�   ��9Eu&9Uu�U�����v����U����A�EtZ�����T��9MuY9UuT�EQQ�$������Y�UY������z���`���u����U����Au��u������E���������؋�^]�����������l$�l$�D$���   5   �   t�������� u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t� ���� ����l$����$����$����l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r �������(��|$�l$�ɛ�l$������l$��Ã�,��?�$�n�����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������,� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����\��Ƀ�u�\$0�|$(���l$�-d������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�L��l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���D��|$�D��<$� �|$$�D$$   �D$(�l$(���D��<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������,� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����\��Ƀ�u�\$0�|$(���l$�-d������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�L��l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���D��|$�D��<$� �|$$�D$$   �D$(�l$(���D��<$�l$$�Q�����0Z�����0Z�������@����������3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u���M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M����p���{L�H��M�����{,�p��2��M�����z�p����M�����z�`���`���������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E�����S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�̔��� "   ]�返��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���x�;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�U�������uV�,���Y�E�^�Ë�|��h��  �u(�  �u�����E ���Ë�U��=p� u(�u�E���\$���\$�E�$�uj�/�����$]�訓��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   �p�3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=p� u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3���L����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-���]���t����-���]�������t
�-���]����t	�������؛�� t���]����jhЛ�_}��3�9��tV�E@tH9��t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�� �e��U�E�������e��U�?}��Ë�U��E��t���8��  uP�O��Y]Ë�U����p�3ŉE�SV3�W��9��u8SS3�GWh��h   S����t�=������xu
���   9]~"�M�EI8t@;�u�����E+�H;E}@�E�������  ;���  ����  �]�9] u��@�E �5�3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w��9  ��;�t� ��  �P��M��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5�SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�,9  ��;�tj���  ���P�M��Y;�t	� ��  �����3�;�tA�u�VW�u��u�u����t"SS9]uSS��u�u�u�VS�u �|�E�V����Y�u������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�8  Y�E���u3��!  ;E ��   SS�MQ�uP�u ��8  ���E�;�tԋ5�SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�8  ��;�t����  ���P��K��Y;�t	� ��  �����3�;�t��u�SW�K�����u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��8  ���u������#u�W����Y��u�u�u�u�u�u����9]�t	�u��+L��Y�E�;�t9EtP�L��Y�ƍe�_^[�M�3��F���Ë�U����u�M��V���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ�p�3ŉE����SV3�W��;�u:�E�P3�FVh��V����t�5���4���xu
jX�����������   ;���   ����   �]�9]u��@�E�5�3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�/6  ��;�t� ��  �P�J��Y;�t	� ��  ���؅�ti�?Pj S�+I����WS�u�uj�u�օ�t�uPS�u���E�S������E�Y�u3�9]u��@�E9]u��@�E�u��5  Y���u3��G;EtSS�MQ�uP�u��5  ����;�t܉u�u�u�u�u�u����;�tV�J��Y�Ǎe�_^[�M�3��D���Ë�U����u�M��T���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v�I���v�I���v�I���v�I���v�I���v�I���6�zI���v �rI���v$�jI���v(�bI���v,�ZI���v0�RI���v4�JI���v�BI���v8�:I���v<�2I����@�v@�'I���vD�I���vH�I���vL�I���vP�I���vT��H���vX��H���v\��H���v`��H���vd��H���vh��H���vl��H���vp��H���vt�H���vx�H���v|�H����@���   �H�����   �H�����   �H�����   �H�����   �uH�����   �jH�����   �_H�����   �TH�����   �IH�����   �>H�����   �3H����,^]Ë�U��V�u��t5�;p�tP�H��Y�F;t�tP��G��Y�v;5x�tV��G��Y^]Ë�U��V�u��t~�F;|�tP��G��Y�F;��tP�G��Y�F;��tP�G��Y�F;��tP�G��Y�F;��tP�G��Y�F ;��tP�pG��Y�v$;5��tV�^G��Y^]��������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U���S�u�M��wQ���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�5����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M���P���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5��N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�����+��;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5��N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3����A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�������   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硰�����3�@�   ����e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+����M���Ɂ�   �ً��]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5��N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�����+��;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5��N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3����A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�������   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�������3�@�   ����e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+����M���Ɂ�   �ً��]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�p�3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u�x{��SSSSS�    ������3��O  �U�U��< t<	t<
t<uB��0�B���/  �$����Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�q%  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �#  =�����/  � ���`�E�;���  }�ع���E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9U�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �;����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�/���Å���/�b�������N�9�����\�U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ë�U���t�p�3ŉE�S�]VW�u�}�f��E��U�� �  #��E��A�#�f�}� �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   t�C-��C �u�}�f��u1��u-��u)3�f9M�f�����$ �C�C�C0�C 3�@�  f;���   3�@f��   �;�u��t��   @uhԔ�Sf�}� t��   �u��u;h̔�;�u0��u,hĔ�CjP������3���tVVVVV艞�����C�*h���CjP�צ����3���tVVVVV�]������C3��s  �ʋ�i�M  �������Ck�M��������3���f�M� ��ۃ�`�E�f�U�u�}�M�����  }����ۃ�`�E�����  �E�T�˃������h  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��z����M�����?  ��  f;���  �]��E�3��ɉU��U��U�U��U�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��U���3�3�f9u���H%   � ���E��[���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �_�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�$���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95����  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�Ë�U��QQ�EV�u�E��EWV�E��  ���Y;�u��e��� 	   �ǋ��J�u�M�Q�u�P���E�;�u���t	P��e��Y�ϋ������������D0� ��E��U�_^��jh��R������u܉u��E���u�ne���  �Se��� 	   �Ƌ���   3�;�|;��r!�De���8�*e��� 	   WWWWW蓒�����ȋ���������������L1��u&�e���8��d��� 	   WWWWW�R�����������[P�j  Y�}���D0t�u�u�u�u�������E܉U���d��� 	   �d���8�M���M���E������   �E܋U��UQ����u�  YË�U���  ��  �p�3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�1d���0�d��VVVVV�    耑��������  SW�}�����4��������ǊX$�����(�����'�����t��u0�M����u&��c��3��0�c��VVVVV�    �������C  �@ tjj j �u�~������u�i  Y����  ��D���  �F?���@l3�9H�������P��4�� ��������`  3�9� ���t���P  ����4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�E���Y��t:��4���+�M3�@;���  j��@���SP��  �������  C��D����jS��@���P�  �������  3�PPj�M�Qj��@���QP�����C��D����|�����\  j ��<���PV�E�P��(���� �4�����)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4������  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@����  Yf;�@����h  ��8����� ��� t)jXP��@����~  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4�����B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4�����b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �|��;���   j ��,���P��+�P��5����P��(���� �4����t�,���;������@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0����t��,�����@��� ��8�������@�����8��� ul��@��� t-j^9�@���u�]��� 	   �]���0�?��@����]��Y�1��(�����D@t��4����8u3��$�_]���    �g]���  ������8���+�0���_[�M�3�^�7����jh���I���E���u�+]���  �]��� 	   ����   3�;�|;��r!�]���8��\��� 	   WWWWW�Q������ɋ���������������L1��t�P�N  Y�}���D0t�u�u�u�.������E���\��� 	   �\���8�M���E������	   �E��FI����u�  YË�U�����h   �p;��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u��[��� 	   3�]�V3�;�|;��r��[��VVVVV� 	   �E�����3���ȃ����������D��@^]ø��á��Vj^��u�   �;�}�ƣ��jP��:��YY�����ujV�5����:��YY�����ujX^�3ҹ��������� ����`�|�j�^3ҹ��W������������������t;�t��u�1�� B��P�|�_3�^��  �=P� t�v  �5���C��YË�U��V�u���;�r"��@�w��+�����Q�M���N �  Y�
�� V��^]Ë�U��E��}��P�]M���E�H �  Y]ËE�� P��]Ë�U��E���;�r=@�w�`���+�����P�:L��Y]Ã� P��]Ë�U��M���E}�`�����Q�L��Y]Ã� P��]Ë�U��EV3�;�u��Y��VVVVV�    �H����������@^]áp���3�9������Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�iY��j^SSSSS�0�ӆ�������V�u�M��#���E�9X��   f�E��   f;�v6;�t;�vWSV�������Y��� *   �Y��� 8]�t�M��ap�_^[��;�t2;�w,��X��j"^SSSSS�0�U�����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�|;�t9]�^����M;�t������z�D���;��g���;��_���WSV�$�����O�����U��j �u�u�u�u�|�����]����������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ��U��j
j �u�'  ��]���U��SVWUj j h���u�*  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    �p�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ�`��SQ�`��L$�K�C�kUQPXY]Y[� ��Ë�U��E��  ��#�f;�u-�EQQ�$�H���HYYtHtHt3�@]�j�jX]ø   ]�% �  ��f��u�E�� u�} t��������]����]����D��z��������@]����%���   ]����������Q�L$+ȃ����Y�  Q�L$+ȃ����Y�  ��U����p�3ŉE�j�E�Ph  �u�E� ����u����
�E�P����Y�M�3������Ë�U���4�p�3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5��M�QP�֋���t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u�脈����YF;�~[�����wS�D6=   w/�������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P���Y;�t	� ��  ���E���}�9}�t؍6PW�u������V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�|��t`�]��[�|9}�uWWWWV�u�W�u�Ӌ�;�t<Vj��2��YY�E�;�t+WWVPV�u�W�u��;�u�u�����Y�}���}��t�MЉ�u������Y�E��e�_^[�M�3��0���Ë�U����p�3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�b���Ë�U��MS3�;�VW|[;��sS������<����������@t5�8�t0�=��u+�tItIuSj��Sj��Sj������3����P��� 	   ��P������_^[]Ë�U��E���u��P���  �P��� 	   ���]�V3�;�|";��s�ȃ�����������@u$�P���0�|P��VVVVV� 	   ��}��������� ^]�jh0���<���}����������4����E�   3�9^u6j
�
C��Y�]�9^uh�  �FP贞��YY��u�]��F�E������0   9]�t�������������D8P���E��<���3ۋ}j
��A��YË�U��E�ȃ����������DP��]Ë�U����p�3ŉE�V3�95��tO�=T��u��  �T����u���  �pV�M�Qj�MQP���ug�=��u����xuω5��VVj�E�Pj�EPV�P�|�T����t�V�U�RP�E�PQ� ��t�f�E�M�3�^���������   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M������E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�����E�u�M;��   r 8^t���   8]��e����M��ap��Y�����M��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�����:���뺋�U��j �u�u�u�������]����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��jhP���9��3ۉ]�j�3@��Y�]�j_�}�;=��}W��������9tD� �@�tP�q  Y���t�E��|(������ P�h����4�c��Y����G��E������	   �E��9���j��>��YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV����YP�]�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�9���P��  Y��Y��3�^]�jhp��8��3��}�}�j��>��Y�}�3��u�;5����   �����98t^� �@�tVPV�>���YY3�B�U�������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��uࡀ��4�V�G���YY��E������   �}�E�t�E��/8���j�J=��Y�j����YË�U���VW�u�M��Y���E�u3�;�t�0;�u,�
K��WWWWW�    �sx�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�[����M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&�iI���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9�uh��P������]����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h���T�áT�V�5���t���tP�֡P����t���tP��^Ë�U��SV�uW3����;�u�H��WWWWW�    �vu������B�F�t7V�!���V����  V�����P�   ����}�����F;�t
P�-��Y�~�~��_^[]�jh���D4���M��3��u3�;���;�u�G���    WWWWW��t���������F@t�~�E��G4���V����Y�}�V�*���Y�E��E������   �ՋuV�����Y�jh����3���E���u�G��� 	   ����   3�;�|;��r��F��� 	   SSSSS�bt�����Ћ����<�����������L��t�P�_���Y�]���Dt1�u�����YP���u��E���]�9]�t�F���M��{F��� 	   �M���E������	   �E��C3����u����YË�U��V�uWV�l���Y���tP�����u	���   u��u�@Dtj�A���j���8���YY;�tV�,���YP���u
����3�V����������������Y�D0 ��tW��E��Y����3�_^]�jh؜�K2���E���u�E���  �E��� 	   ����   3�;�|;��r!�E���8�mE��� 	   WWWWW��r�����ɋ���������������L1��t�P�����Y�}���D0t�u�����Y�E���E��� 	   �M���E������	   �E���1����u�,���YË�U��V�u�F��t�t�v�=���f����3�Y��F�F^]�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%�������������h� ���Y����̃=l� uK�d���t�`��Q<P�B�Ѓ��d�    �p���tV���@6��V�*r�����p�    ^�                                                                                                                                                                                           8� N� `� l� |� �� �� ��  ֞ � � $� 8� F� R� `� j� �� �� �� �� �� ҟ � � � � 0� J� b� |� �� �� �� Ƞ ֠ �  � � 0� <� T� l� |� �� �� �� �� �� ʡ ֡ � �  � 2� B� X� h� z� �� �� �� �� Т � �� � � "�         �         �63E�m�        `���                    ۪�O       w   Е �{ bad allocation  *** (c)2012 Michael Auerswald   There was a problem registering the Point Position plugin.  *** Point Position v0.3 *** C4DSDK - Edit Image Hook:   -SDK is here :-)   -plugincrash    -SDK executed:-)   -SDK    -help   --help  c:\program files\maxon\cinema 4d r13\resource\_api\c4d_general.h              �c:\program files\maxon\cinema 4d r13\plugins\pointposition\source\pointposition.cpp     �� �k �k  l l  l �k 0l Pl `l @l �l �l �l �l pl �l � � � � @� P� �  � `� p� �� �� �� � �  � �  � 0� @� PointPosition   VPpointposition %s     c:\program files\maxon\cinema 4d r13\resource\_api\c4d_file.cpp c:\program files\maxon\cinema 4d r13\resource\_api\c4d_resource.cpp #   M_EDITOR    D��k res -DT�!��-DT�!�?      �?-DT�!	@        -DT�!@�h㈵��>{�G�zt?      �?       @      �A      �A
ףp=
�?       �
ףp=
�?      @      @����MbP?c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basebitmap.cpp   X� � c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gv\ge_mtools.cpp ԗP� ��� h��� �� 3� 3� ����                   �?      �?3      3            �      0C       �       ��              e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    ��@�EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                                              �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �      �?5�h!���>@�������             ��      �@      �                                                  �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������              �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC              ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=      �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow       8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �              8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7�������             ��      �@      �        	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =   ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx           Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        �p�p�p�p�p�p�p�p�p�p�j�k�k�k�klk�p�p�j�p|pxptppplp`p\pXpTpPpLpHpDp@p<p8p4p0p,p(p$p pppppppp p�o�o�o�o�o�o�o�o�o�o�o�o�o�o`o@o o o�n�n�n|n\n4nnnn�m�m�m�m�m�m�mhm@mm�l�l�l�l`l4ll�k�jGetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL     �U��?�wB%�K�=      �?   �[��?(�6N�g�=      �?   $�?V�`t� >      �?   ��տ?��2n{a>      �?   ����?��M��=      �?   H{��?{4�r>      �?   Pא�?"�"�>      �?   �u[�?��*��>      �?   ����?G�0��_(>      �?   4wb�?��i^^?(>      �?   ��0�?p3���>      �?   @��?F��M>      �?   8M��?�B�V��>      �?   ��d�?}B��a.>      �?   ȴ�?d�����>      �?   g��?�ߊ��>      �?   �@�?�f\���*>      �?   �~e�?�-��f>      �?   �]%�?D	�G��?>      �?   ���?�\����>>      �?   X���?�1��#>      �?   �E�?��h��>      �?   �?��?�ⳇ��>      �?   ����?�$	�49>      �?   x�8�?k���0H<>      �?   ����?r��ش8>      �?   8fm�?�"m>">      �?   ħ �?[��<c�'>      �?   �k��?"���%>      �?   ���?݉@fR�8>      �?   ����?��T���:>      �?   T�!�?3&�F>      �?   � ��?<����[#>     ��?   �%�?�Y:/(A6>      �?   ����?��N��2>     ��?   8O�?�r�!'	>      �?   ��r�?���8{K>     ��?   �p��?9��l�9$>      �?   �
G�?�aj	�i9>     ��?   T|��?'\�|#<>      �?   $��?�}�dj�#>     ��?   �Wn�?׈MVx:>      �?   ,���?1�8o,>     ��?   D�$�?	c�/�
>      �?   @ |�?��x7|�1>     ��?   |���?��9>      �?   p #�?�IA��u=>     ��?   �s�?�x ٴ4>      �?   p���?edf�&�.>     ��?   ,�?��f���A>      �?   h�*�?v����2>     ��?   $gN�?RE\��K>      �?   �q�?'^��IE>     ��?   DΒ�?��&a��H>      �?   L���?�&KrQF>     ��?   ,���?�#/�'�>      �?   إ��?]X�c�?>     ��?    ��?�Ԯ}�>      �?   �e.�?�IdW�A>     ��?   �K�?���ΐ?>      �?   Xg�?��4*�A>     ��?   _��?�[�ǆJ>      �?   ���?1���0H>     ��?   ���?�hc#�]G>       @   ,*��?�Q�x
�F>     @ @   p���?ek�R�.N>     � @   �� �?�Ӿ�n@>     � @   �b�?�����O>      @   $Q/�?CJ���O>     @@   ��E�?������G>     �@   �[�?�3E�{A>     �@   T�p�?�SfI�S:>      @   X΅�?B6)�1�<>     @@   �3��?>ځ���7>     �@   $��?s(��N>     �@   @���?V�
6�f=>      @   (���?��{��>     @@   (W��?��-�Jg >     �@   ����?��"a�PK>     �@   xm�?,S��ڤ6>      @   ���?�6��hb">     @@    �-�?�k,�<>     �@   X�>�?�0����=>     �@   �O�?�׀IX�H>      @   �-_�?���
@>     @@   ��n�?���2E>     �@   �P~�?�=�ő�8>     �@   lj��?�[j&,>      @   L7��?��x��82>     @@   ����?c�#V�B>     �@   0��?7ڨ.�Y>     �@   P���?�[�p&>      @   ؔ��?h4�M��A>     @@   � ��?E�p�l E>     �@   �+��?�o�$�E>     �@   h��?\���*�K>      @   ���?-�?��B>     @@   P8�?�(l�|�@>     �@   �p!�?u���@�J>     �@   @p-�?�V��1>      	@   �89�?����5>     @	@   <�D�?��ƀ�7>     �	@   h)P�?R`D�OG>     �	@   �T[�?9%� ��K>      
@   �Mf�?��/�<>     @
@   �q�?�Ò��?>     �
@   �{�?4��2G<>     �
@   L��?Â���|/>      @   �Y��?���s�
@>     @@   �k��?��Ò�a@>     �@   XS��?x(3��u8>     �@   ���?v�O,ib>      @   ȥ��?�&L͒C>     @@   ���?��}��L>     �@   �X��?Lo����>     �@   �x��?-�Ϡ�9>      @   �s��?6FID?9>     @@   8J��?����gsL>     �@   d���?��y>     �@   ���?>�&�09C>      @   ����?
��<�A>     @@   (J�?I�V	C>     �@   `w�?��^@�N>     �@   ���?�#��%�@>      @   �s�? �M�K>     @@    D'�?ή�Q��->     �@   ��.�?9!���G>     �@   ��6�?.����1>      @   >�?.1�NcB>      @   �cE�?�sǔ�1>     @@   L�L�?�n�HN>     `@   H�S�?�W��$>     �@   8�Z�?
Ȃ�q�;>     �@   ��a�?N�/�[7>     �@   (�h�?�=�mC>     �@   0oo�?�H75M>      @   Hv�?P��.�#>      @   �|�?�G���7>     @@   �*��?�#4��2I>     `@   ����?o���oJ>     �@   ����?���-��#>     �@   ���?�h��%F>     �@   @��?R�x^D>     �@   PP��?�� s�@>      @   4L��?P�_!
�#>      @   4��?��:#�G>     @@   L��?qg�:&J>     `@   Hɹ�?5L$.��4>     �@   \w��?!�1�C>     �@   ���?���[<>     �@   D���?��<���=     �@   ���?��
~���=      @   �y��?������B>      @   ����?�~.���4>     @@   h��?��u�|�8>     `@   �E��?A8yL;>     �@   �h��?��41��C>     �@   �{��?-���+oF>     �@   $��?x���O>     �@   s��?�՝m�T2>      @   �W��?����=>      @   �-�?î�\�=>     @@   ��?���\=�=     `@   ��?j\&">     �@   �X�?��1�D>>     �@   ���?�#O#`�I>     �@   ��?�}���0>     �@   ��?���F\IE>      @   t{#�?��ׯ,B>      @   0�'�?�E� ]�$>     @@   ,>,�?��ކ?5>     `@   ��0�?��iIqE>     �@   ��4�?�ha�;>     �@   �9�?��A���D>     �@   �.=�?̤KF�w�=     �@   DMA�?�����=      @   `E�?ap�I0�H>      @   �gI�?��:���->     @@   �cM�?��%Q>     `@   @UQ�?Ly5ښoE>     �@   �;U�?v�g�0�/>     �@   �Y�?jv�U�G>     �@   �\�?�����yK>     �@   ,�`�?A%My��>      @   md�?���H>      @    h�?�p���M>     @@   0�k�?k��}<>     `@   �ho�?����f7O>     �@   ��r�?���}�O>     �@    �v�?+��i�I>     �@   @z�?�b�B'=>>     �@   `�}�?Z����M>      @   ����?1�����M>      @   �a��?R�~���=     @@   t���?QNT	��B>     `@   x��?�W3c�L>     �@   g��?�+(����=     �@   D���?q���J�K>     �@   L��?� ;,*>     �@   8!��?������D>      @   ,O��?� ����E>      @   Du��?��in]D>     @@   ����?%����3F>     `@   P���?^��F"VM>     �@   ����?�}�30}->     �@   @���?�~F	y�;>     �@   ����?l	R(>     �@   躰�?��\�7`>      @    ���?�dg���;>      @   ���?�;Sv�@E>     @@   <|��?�����M>     `@   �Y��?|}�;�2>     �@   ,0��?�<v��G>     �@   $ ��?̯�/p�">     �@   ����?���\(0>     �@   |���?[s$���F>      @   I��?�d�ӔV>      @   T���?���0)LK>     @@   h���?�)�5G�5>     `@   XY��?�|��zJ>     �@   @���?W�޾�L?>     �@   0���?����6:>     �@   <3��?��Q���B>     �@   x���?7o��/�M>      @   �Q��?�Kc�Z�0>      @   ����?�z-�A5>     @@   Z��?"B�DcI>     `@   ����?��`I�.>     �@    L��?L�d�%>     �@   ���?"�l"w �=     �@   �(��?�?��!>     �@   ���?��j^�J>      @   8���? ϞH��0>      @   LL��?���%�C>     @@   T���?��J�+N>     `@   d���?;l�>�0>     �@   �B��?�^{v�@>     �@   Ȋ��?�@Y˕B>     �@   @� �?T�l���0>     �@   ��?w4n4>      @    G�?�oN�=�;>      @   h|�?�L�{�/>     @@   <�	�?B�nu5>     `@   ���?���`�,+>     �@   d�?����5>     �@   �$�?l��  >     �@   �C�?~+^��M>     �@   �^�?�PK�QD >      @   ,u�?^{�#tF>      @   |��?�^4K�� >     @@   ���?��4�O
>>     `@   ���?XEړ� J>     �@   ���?(�gԹ�,>     �@   �� �?43-spF>     �@   ��"�?P`E5�+*>     �@   ��$�?=�QQ�D>       @-DT�!�?\3&��<_nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                                                                                                                                                                                                                                                                                              ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           p� �   RSDSNI�A�B�V�7 Y�d   C:\Program Files\MAXON\CINEMA 4D R13\plugins\pointposition\obj\pointposition_Win32_Release.pdb             X�d���    �       ����    @   H� �        ����    @   ��           ����               ĖԖd���    8�       ����    @   ��            T��           �(�Ԗd���    T�       ����    @   �             ���            ��l�           |���    ��        ����    @   l�           ����    ܰ        ����    @   ��            ���           �� �    ��        ����    @   �            �0�           @�L���    �       ����    @   0�            @�|�           ����    @�        ����    @   |�            |�Ę           Ԙܘ    |�        ����    @   Ę        �1 �� ��                     ����    ����    �����     ����    ����    ����    f    ����    ����    ����    P    ����    ����    ����    y    ����    ����    ����    =    ����    ����    ����     ����     ����    ����    ����    �!����    �!����    ����    ����    J'    ����    ����    ����**    ����    ����    ����    d4    ����    ����    ����x5�5    ����    ����    ����    �7    ����    ����    ����    �i    ����    ����    ����    ym    ����    ����    ����    �p    ����    ����    ����    J�    ����    ����    ����    ��    ����    ����    ��������    ����    ����    �������    ����    ����    ����    ��    ����    ����    ����x���    ����    ����    �����2�    ����    ����    ����    E�    ����    ����    ����    T�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    k�        7�����    ����    ����    u�    ����    ����    ����    W�    ����    ����    ����    ���         6�                       8� N� `� l� |� �� �� ��  ֞ � � $� 8� F� R� `� j� �� �� �� �� �� ҟ � � � � 0� J� b� |� �� �� �� Ƞ ֠ �  � � 0� <� T� l� |� �� �� �� �� �� ʡ ֡ � �  � 2� B� X� h� z� �� �� �� �� Т � �� � � "�     �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �GetLastError  �HeapFree   GetProcAddress  �GetModuleHandleA  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �InterlockedIncrement  �SetLastError  �InterlockedDecrement  !Sleep ExitProcess �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA � DeleteCriticalSection �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW zWideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  �LeaveCriticalSection  � EnterCriticalSection  TVirtualAlloc  �HeapReAlloc �WriteFile [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �RtlUnwind �LoadLibraryA  �InitializeCriticalSectionAndSpinCount ZRaiseException  �GetLocaleInfoA  �LCMapStringA  MultiByteToWideChar �LCMapStringW  =GetStringTypeA  @GetStringTypeW  �SetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW x CreateFileA C CloseHandle AFlushFileBuffers  KERNEL32.dll                  ۪�O    ��          x� |� �� �  ��   pointposition.cdl c4d_main                                                                                                    ||    .?AVNodeData@@      .?AVBaseData@@      .?AVVideoPostData@@     .?AVPointPositionPostData@@ ||||||||||||||||||    .?AVGeToolNode2D@@      .?AVGeSortAndSearch@@       .?AVGeToolDynArray@@        .?AVGeToolDynArraySort@@        .?AVGeToolList2D@@  |||u�  s�  N�@���D|    .?AVtype_info@@             sin             cos             atan            log             sqrt            asin            acos            �|�|�|�|�|�|�|�|�|�||    ��������b'    �����
                                                                   x   
                                                                                                                                                                                                                                                                                            �   �	   �
       �   �   �   T      �   �   �   \   <   �    �!   �"   x   �y   �z   ��   ��   �                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                        ���5�h!����?      �?             ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          R-H2HAS  ?  atan2        |b�b_H�b�b�b_H�b]H]H�H]H�b�b_H�H                                                                                                                                                                                                                                                                                                                                                   abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ������C                                                                                              �            �            �            �            �                              p�        ��������   ��        k�j               
      p?  �?   _       
          �?      �C      �;      �?      �?      ���������������������ΞӞ��
��.�>�^�c�}�������Ο���!�&�F�Z�r�������Šʠ����*�J�O�i�n�������Ρ����2�F�^�r���������֢��  �&         8:   <:   ,:   0:   x�   p�!   h�   $:   :   :   `�   X�   �9   �9    �9   :   �9   P�   �9   H�   @�   8�   0�   (�"   $�#    �$   �%   �&   �      �      ���������              �       �D        � 0     ����    ��������������������|�p�h�\�X�T�P�L�H�D�@�<�8�4�0�,�$����H� �����ܓГē����������	         ��.   l�������������������p�   .         ���5      @   �  �   ����             ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �            �p     ����    PST                                                             PDT                                                             ��������        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
   ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l          ��������                                                                                                                                                                           �   0040E0t0�0�0�0�0�0�0�01#151G1a1s1�1�1�1�1�1�172x2�2�23,3E3�3�3�3�3�3)4;4L4t4�4�4�4�4
5=5K5^5s5�56'6Y6y6�6�6�6�6*7�7�78�8
99%969H9Z9q9�9�9�9:':4:Q:d:�:�:�:;!;D;d;�;�;�;<D<t<�<�<�<=$=D=d=�=�=�=�=�=>!>1>D>d>�>�>�>??$?d?�?�?�?�?      �   0010A0T0t0�0�0�0�01?1d1�1�1�1�1�1242_2�2�2�23*3T3t3�3�3�3�3444T4t4�4�4�445t5�5�546t6�6�6�6!7A7T7�7�7�7�7�78$8D8d8�8�8�8"9H9e9�9�9�9�94:R:f:v:�:�:�:�:;4;T;t;�;�;�;�;<$<]<r<�<�<�<�<=#=D=^=r=�=�=�=�=�=>(>A>o>�>�>�>??'?6?d?|?�?�?�?�?   0    040]0�0�0�0�0+1>1t1�1�1�12$2D2d2�2�2�2�2�23$3d3�3�3�3�34$4D4d4�4�4�4�4�45!545d5�5�5�5�5�5�56&686T6�6�6�6�6�6�67747E7S7q7�7�7�7�78848L8`8p8�8�8�8�8�8�8949L9`9o99�9�9�9::$:D:d:�:�:�:�:�:;$;T;t;�;�;�;�;<A<T<�<�<�<�<�<=4=Q=a=q=�=�=�=�=>$>D>d>�>�>�>�>�>?D?^?u?   @     g0�0�0�0�0�0�0�1�1�1�12D2d2�2�2�2�23$3D3a3t3�3�3�3�3414D4_4m4{4�4�4�4�4�4 5!5D5d5�5�5�5�5�5�5�56/6=6K6Z6l6�6�6�6�6747T7t7�7�7�7 88-8W8i8�8�8�8�8�8949T9t9�9�9�9�9�9�9:4:N:b:q:�:�:�:�:�:;,;=;K;b;w;�;�;�;�;�;<<&<t<�<�<�<�<=4=A=Q=d=�=�=�=�=>$>D>d>�>�>�>�>?$?D?d?�?�?�?�? P     0$0D0d0�0�0�01$1D1d1�1�1�1�12$2D2d2�2�2�2�23$3D3d3�3�3�3�34$4D4a4t4�4�4�4�45!515A5T5t5�5�5�5�56$6I6j6�6�6�6�7�788-8`8u8�8�89(979k9�9�9�9+:f:�:�:�:�:�:�:;;&;9;K;];o;x;�;�;�;�;�;<%<8<d<r<<�<�<�<�<�<�<=$=6=R=h=�=�=�=�=�=�=>">3>F>t>�>�>�>�>�>�>�>�>?4?F?b?x?�?�?�?�?�? `  �    0020D0V0_0}0�0�0�011171I1[1m11�1�1�1�1�12$262H2Q2o2�2�2�2�2�2�23.3D3b3o3�3�3�3�3�34D4a4�4�4�455 5;5W5p5�5�5�5�5666X6u6�6�677$7}7�7�7�7�7�7828O8�8�849I9k9�9::1:A:T:�:�:�:�:�:;4;Q;d;�;�;�<==�= >'>.>5><>C>J>Q>X>_>f>m>t>{>�>�>�> p  �   /0Q0|0�0�0�0S1e1�1�1I2e2�2�2I3l3�3�3�3�34%4�4�4!5|5�56$6D6d6�6�6�6�6�9�9�9G:O:h:�:�;�;�;�;�;�;�;�;<><�<�<=A=�=�=Q>�>�>K?�?   �  �   0F0W0�0�0�0�0�01b1s1�1�1�1�1�1�1 2�2\6`6d6h6l6p697P7a7P8�8�9�9�9�9�9::5:_:�:�:�:�:�:;;5;_;�;�;�;�<�<	==&=i=�=�=8><>@>D>H>�>?1?D?q?�?�?�? �  �   40d0�0�01$1D1a1�1�1�12$2Y23$3D3{3�3�3	4$4�4�4�4+5^5y5�5�5�56$6T6t6�6�6�6747F7t7�7�7�7�8�8959u9�9�95:�:�:�:;E;�;�;<M<�<�<=R=�=�=>E>�>�>?R?�?�?�?   �  �   20e0�0�051u1�1�182S2�2�2�2�23U3�3�34e4�4�4A5i5�5�5�5�5�56B6j6�6�6�67X77�7�7"8e8�8�8�89R9�9�9�98:v:T<�<�<�<�<�<�<=====$=+=2=9=@=G=N=U=\=�>�>�>??3?:?T?n?�?�?�?�?�?�?�?�?�?   �  �   0!0D0a0�0�0�0!141a1�1�1�1�1232F2q2�2�2�23$3T3�3�3�3�3�3$4d4�4�4�4�445T5q5�5�5�5�56D6v6�6�617D7t7�7�7�7�9
::@:;&;�<�<�<$=T=t=�=�=�=�=�=>4>d>�>�>�>�>�>!?D?a?�?�?�?�?   �  �   0�0,1�1�1�1�2�2�2�3�3�34Q4[4�4�45$5Q5t5�5�5�5�5646a6t6�6�67!7A7a7�7�7�7818Q8t8�8�89!9D9d9�9�9�9�9:$:D:d:�:�:�:�:�:;4;�;�;�;L<w<�<�<Q=�=�=>�>�>�>A?^?v?�?   �  �   0#0�0�0�0!1D1�132\2�23,3T3�3�3$4�4�4�4K5�5�5A6g6�6�6A7g7�7,8�8�8�8n9�9�9:>:S:�:�:;|;�;<4<Q<a<t<�<�<�<=$=T=t=�=�=�=>4>Q>t>�>�>? ?B?~?�?�?�?   �  �   00Q0q0�0�0�0�0�1�1�1�1�1�1242Q2d2�2�2�2�23D3t3�3�3�3�3�3444W4�4�4�4'5b5�5�5�6�6�6D7t7�7�7�;=<M<|=�=>D>K>f>�>�>�>?]?�? �  �   0'0D0d0�0�0�0�011$1A1Q1d1�1�1�1�1�1242T2x2�2�2�2�2$3D3d3�3�3�3�34$4d4�4�4�4�4�455A5_5�5�5�5�5646T6�6�6�6�6�67!747T7i7}75>:>@>D>J>N>T>X>^>b>g>m>q>w>{>�>�>�>�>�>�>�>/?4?>?r?�?�?�?�?�?�?   �   /0K0c0�0�0P1[1�1�12232�233o3u3�3�3�3&484�4�4�4�45i5w5�5�5�5�5�5�526�6�6�6�6�6�67"7b7�7�7�788/8B8�8�899D9h9s9�9�9�9":-:?:R:�:�:7;Q;Z;b;�;�;C<U<{<�<�<�<�<=�=�=�=�=>!>+>B>^>??2?=?    �   �1d2�2�7�8U:�:�:�:�:�:�:�;�;�;�;�;�;<<<<<$<+<3<;<C<O<X<]<c<m<v<�<�<�<�<�<�<�<�<�<�<�<�<�=�=�=�=>>->4>[>a>l>x>�>�>�>�>�>�>�>�>�>�>???#?/?5?B?L?S?k?z?�?�?�?�?�?   \  ,020\0b0~0�0�061Y1c1�1�1�1�1222'2-2B2P2[2b2}2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 333*353:3E3J3U3Z3g3u3{3�3�3�3�3�344I4R4^4�4�4�4�4�45!5'50575Y5�5�5�5�5�5�5�5666.696S6_6g6w6�6�6�6777767�7�7�7�788E8�8�8�8�89/9p9�9�9:
:.:L:n:y:�:�:�:;%;/;@;K;�<==="=(=�=�=�=�=�=�=�=�=)>x>�>�>�>�>�>??D?I?W?_?k?r?{?�?�?�?�?�?�?�?�?�? 0 �   e0k0�0�0U1r1�1�2�2�2�2+3E3h3u3�3�3�3�3�3�3�34P4V4^56!6(626\6j6p6�6�6�6�6�6�6�67�7�7�7�7:&:,:F:K:Z:c:p:{:�:�:�:�:�:�:�:�:�:�:�: ;;;;+;2;8;F;M;R;[;h;n;�;�;�;�;<�?�?�? @ �   0P0�0h2s2{2�2�2�2�2"3+323;3{3�3�3�3�344/4S4~4�4�4�45555@5�5�5�5�5�5�5�56S6_6�6�6 7I7�7X8�8+9,:<:M:U:e:v:;%;5;A;^;d;y;�;�;�;n<�<�<�<�<�<
=="=N=l=x=�=�=�=�=�=�=�=�=>'>;>V>g>p>�>�>�>�>�>�>�>???/?F?M?�?�?�?�?�?�? P �   Y0e0y0�0�0�01171G1S1b1$2n2�2�2353I3T3�3'4/4<4�4�4	55-595E5Q5v55�5�5�5�5�5�5�5�56
66"6+646s6w6{66�6�6�6�6�6�6�6�6�6�67�7�7�78!8M8U8x8�8�859A9a9q9}9�9�9::~:�:�:�:;
;;G;v<~<�<"=*=6=�=�=�=�=�=>�>�>�> ???�?�?�?�? ` �   70?0G0S0_0�0�0�1�1!2)2�2$3a3�3q4�4�4�4�4�4�5�5�5�6�6�6O7�7�79'9a9n9x9�9�9�9�9�9�9�9::<:s:�:�:+;H;�;�;<�<�<�<�<�<�<�<==8=A=G=P=U=d=�=�=�=�=�>�>"?n?�?   p �   0k0�0�0�0�01�1�1�12232�2�2�34�4�5�5�5�5�5�5 66-6S6q6x6|6�6�6�6�6�6�6�6�6�6�6�6V7a7|7�7�7�7�7�7�78888 8$8(8,808z8�8�8�8�8S;X>_>j?   � `   0*0P0�0�0�0)45�6�6�6�8�:�:�:�:�:�:�:�:�:;!;-<V<�<�<===t=�=�=J>P>�>�>�>�>"?(?4?{?   � �   (0-0?0]0q0w0�01"10151:1?1O1~1�1�1�12"2)2.252:2�2�2�2B3Q3Z3o3�3Z4�4�4�4�4�4�4�4�451585<5@5D5H5L5P5T5�5�5�5�5�56!6<6C6H6L6P6q6�6�6�6�6�6�6�6�6�6�6:7@7D7H7L7�7�7�7�7�7�7�78888*838B8G8Q8_8�8�8�8A:H:N:�:�;�;Y<�<�<=?=�=�=�=�=�=X>�>   � 4   �5�6�657�7�78=8�9�9�9�:�:�:=z>�>�>�>�>4?   � l   =0�0�0C1�1�3�3�3�3�3474�4�4�4�4�4�4�4�4,5�5s6�67�7m8w8�8�8�8�8�8�8�8�9�9<<+<M<_<q<�<�<�<�<�>�?�? � T   �0r122�2�2�2i3�3#45!5�5�6O7U7�7�78�8�8�8�9Q<h<�?�?�?�?�?�?�?�?�?�?�?�?   � $   V102J2Y2�2�2	3=�>??9?w?�? � x   _0�0x1�1�2�2
3�4x5A6r6�6�6�6�7�7�7e8�8�899,9;9H9T9d9k9z9�9�9�9�9�9�9�9:O:^:g:�:�:�:�:)<G<�=�=	>�>�>�>�?�?�?   � �   0$011�1j3z3�3�344W4s4�4�455$525:5G5e5o5x5�5�5�5�5�5�5{6�6N7o7{7�7�7�7�7�8�8�8�8=9�;�;P<V<[<a<h<z<=�=�=�=>>x>�>�>�> ?4?c?        �0�0�0�011 1;1  �    1,1014181<1H1L133 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3l4p4�5�5�5�5�5�5�5�5 66666�6�6   p �   111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2 � �   �5�5T6X6\6d6|6�6�6�6�6�6�6�6�6�6�6�6 77777 7(7@7P7T7d7h7x7|7�7�7�7�7�7�7�7�7�7�7 88(8,8<8@8D8L8d8t8x8�8�8�8�8�8�8�8�8�8�84989X9x9�9�9�9�9 ::(:D:H:h:�:�:�:�:�:;(;H;d;h;�;�;�;�;�;�;�;<(<H<h<�<�<�<�<�<   � �   000 080T0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01@1\1`1d1x1|12222 2$2(2,2024282H2�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4j6n6r6v6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6; <h<x<�<�<�<�<�<�<�<�<�<�<�< ==n=r=v=z=~=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>
>>>>>>">&>*>.>2>6>:>>>B>F>J>N>R>V>Z>^>b>f>j>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � X    00000000 0$0(0,0004080<0@0D0H0L0P0T0X0h0p0t0x0|0�0�0�0�0�0�0�0�0�0 44                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  