MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��<�b�o�b�o�b�ok,o�b�o��o�b�o��5o�b�o�o�b�o�b�o�b�o��4o�b�o��o�b�o��o�b�oRich�b�o                        PE  L /��T        � !
  $  �      �      @                       @    ��  @                   �� \   � (      �                    *  @L                            �� @           �� �                          .text   �#     $                   `.rdata  o   @  p   (             @  @.data   �;   �     �             @  �.idata  )
   �     �             @  �.rsrc   �         �             @  @.reloc  �/     0   �             @  B                                                                                                                                                                                                                                                                                                        ������F5  �!3  �|  �wS  �4  ��  �(G  �35  �  �9
  ��  �?  ��6  �D  ��?  �k  �7  �  �\7  ��  �  �K  ��0  �  �;  ��:  �t5  �5  �
!  �54  �	  �3  �F4  ��6  �<  �'J  �BB  �}#  ��9  �SO  �2  �
  �t<  ��	  ��9  ��  �@>  �N  ��	  ��4  �  �R  �"  �  �G  �C1  �~A  �y  �$:  �6  �j>  ��?  �  ��  �F  ��  �  �g?  �27  ��E  ��9  �  �2  �  ��  �?3  �Z:  ��/  �P  �  �VG  ��4  �I  �3  ��  �5  �8B  �s4  �.K  �  �1  �o3  �  �55  �  �KA  �1  �5  ��9  �wI  �L  �L  �9  �c  �  ��1  ��0  �  �z  ��/  �  �{9  �M  ��  �LC  �;  ��  ��5  �2  �#9  �n  �   �t4  �  �  �53  �@1  �{4  �  �  �  �1  �R  �  ��:  �	  ��.  ��I  ��
  �=  �J  �.  � G  �k  �;  �  �0  ��
  �0  �2  �@  ��0  �  ��0  ��D  �O1  �;  �  �  �k/  �vE  �a  �L	  �W2  �2  �9  �(F  �9  �^/  �Y  �L  ��	  ��  �E1  �p  �  �&G  �Q  �l  �  �b  �]  �A  �#/  �.  ��  ��@  �@  �  �e	  ��
  �  �6/  ��>  ��  �3  ��  ��2  �H:  ��  �n:  �4  �  �?  �Z  ��  �  �  ��  ��  �2  �w  �  �]K  ��=  ��  �?  �YK  ��  ��-  �/  �  �   �.  ��  �  �0  ��  �  ��8  ��K  �9  �  ��  �  ��B  ��8  ��,  � ;  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��W�}OxS�]V�u����uOy�^[_]� �������������������������������������������U��E�� tHt3�]ù����V  �����]ø   ]����������������������U��E�M;�|��]���������������������P�X����U���E����E�X�E�X]� ������U��M��E�E������A���X�I�X]�������������U��M�U���E��A�B�X�A�B�X]�����������U��EE]������U��E#E]������U��EE]������U��E#E]������U��E#E]�����������P�P�P�P �P(�P0�P8�P@�PH�PP�XX�������������������������U��E��E	]������������������U��E]���������U�조�V��H�QV�ҡ���H�U�AVR�Ѓ���^]� ����������������U�조�V��H�QV�ҡ���U�H�E�IRj�PV�у���^]� �������������������������̡���P�BQ��Y����������������̡���P�B<����̡���P�B<�������������������̋��     �@    �����������������U����M�    �H]� �����������U��UV���    �F    ������   �Aj RV�Ѓ���^]� ���������������������������̡�����   �Q��Y���������������U�조����   �E�RPQ�MQ�҃�]� �������������U��E�M�UP���   QR�� ��]������������������U��U��t�M��t�E��tPRQ�`� ��]�����������̡���P�B �����U�조��P�R$]�����������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��E�P�E���   ���$P��]� ������������U�조��P�R0]�����������������U�조��P�R4]�����������������U�조����   �R]��������������U�조����   �R]��������������U�조��PH�EPQ���  �у�]� ����������������̡�����   ���   ���������������U�조����   ���   ]����������̡�����   ���   ���������������U�조����   ���   ]�����������U�조����   ���   ]����������̡�����   ���   ���������������U�조��P|�EP�EPQ�J�у�]� ����������������U�조��P|�EPQ�J�у�]� �������������������̋�������������̡���Pd�Q�Ѓ�����������������U�조��Pd�EPQ�JX�у�]� �������������������̡���Pd�BQ�Ѓ���������������̡���Pd���   Q�Ѓ������������̡���Pd���   Q�Ѓ�������������U�조��Pd�EPQ�J�у�]� ��������������������U�조��Pd�EP�EPQ�J�у�]� ����������������U�조��Pd�EPQ�J`�у�]� ��������������������U�조��Pd�EP�EPQ�Jp�у�]� ����������������U�조��Pd�EP�EP�EPQ���   �у�]� ���������U�조��Pd�EP�EP�EPQ�Jt�у�]� ������������U�조��Pd�EP�EPQ���   �у�]� �������������U�조��Pd�E���   ��VPQ�M�Q�ҋu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у���^��]� ���������������������������U��E����]� ����������������U�조��PH�R,��`VW�E�P�ҋ��E�   ���_^��]� �����������������U�조��PH�EP�EPQ��p  �у�]� �������������U�조��PH�EPQ���   �у�]� ����������������̡���PH���   Q�Ѓ������������̡���PH��p  j h�  Q�Ѓ���������������������̡���PH���   h�  Q�Ѓ�������̡���PH��p  j h�  Q�Ѓ���������������������̡���PH���   h�  Q�Ѓ�������̡�����   �B(������������������U�조��HD�A,]�����������������U�조��HD�A0]����������������̋���������������U�조��H�U���  h�Mj{R�Ѓ�]� �����������U��EP��Q  ��]� ������������̋�� ������������U��E�3�;��]� �������������U���UV�����   W�:3���3��S��z�����   3���3��S��z��%�   3ǋ��S��3Ɖ�R�����   3���3��S_�^]� ���������������������������������������̋�� ������������U��EVP���������^]� ����������U��EVP��������^]� ����������U��E��U3�;
��]�������������U��M�E9s���;�r��]������̋�������������̋A�������������U��E�;u�@;Au	�   ]� 3�]� �������������������A�����������������������U��V�uW�}��MQ�ΉE������W�EP�ΉU�����_��^]���������������U��E���3  SVW�$�( �E�M�U��M�P�U�H�M �P�U$_^�H�P[]ËE�M�U�H�M�P�U�H �M �P$�U$_^�H(�P,[]Ã}( �Et>�M�U�u�}�] �H0�HH�M �P4�PL�p8�pP�x<�xT�X@�]$_�HX^�XD�X\[]ËU�M�P0�U�H4�M�P8�U �H<�M$_^�P@�HD[]Ã}( �E�M�U�HH�PLt2�u�}�] �H0�P4�U �p8�pP�x<�xT�X@�]$_�PX^�XD�X\[]ËM�U�HP�M �PT�U$�HX�P\_^[]��& ' @' �' ��������������������������������������������������������������������������������������������U�조�VW�}��Hd���   Vh�  W�ҡ���Hd���   �VRh�  W�Ћ���Qd���   �� VjW�Ѓ�$_^]� ������������������������������������U��S�]V�uW�}�����Ox��$    +���UOy�_^[]� ���������������U��E���X�@�����@    �     ]����������������U��E�8 t�x |�   ]�3�]�����U��E�P�M;Qu� ;u�   ]�3�]���������������U�조��P�B$V�uW��h�Y ���Ћ���Q�B0jh�  ���Ћ���Q�B4j
h�  ���ЋMVQ���^  _^]� ��U��QSV����ًHH���   h�  S�҉E�����HH��p  j h�  S�҃��؋E�����   ;���   ��xg;�}c����Qd�M���   j �v�u��QPV�E��ҋ���Qd���   ��ËEj PSV�ы���M��Bd�Ptj SQV�҃�0^[��]á���Hd�U���   j R�v�ËERP�у�^[��]Å�x);�}%����Bd�M���   j Q��ӋUQR�Ѓ�^[��]������U���EW���    �    ty�E   tpjW���h  ���t`���t
S�a  ��~D���tJ����QHh�  P���   �Ѓ���~ �����QHh�  P���   �Ѓ����    �    �Et5�> u0����QH���   S�Ѓ���t����QH���   S�Ѓ������   ����QH���   S�Ѓ�����   �> ��   ����QH���   S�Ћ���QH�����   h�  W�Ћ���QH�E���   h�  S�Ѓ�9Eu7����QH���   h�  W�Ћ���QH�����   h�  S�Ѓ�;�t�    _]Ã> u�_]����������������j jP�֛ �����U��V�u���"�  ��t
��t��uz������   ���   ��jP�ΉE��  ������   �M���   �Ѕ�~%������   ���   �EP�у��   @^]� ������   ���   �MQ�҃�3�^]� ��U���   ��3ŉE��ESV�u�ًM�i  �{ �_  �C����R|Wh�  QP�B�Ћ������$  ;{�  ����QH���   h�  W�ЋK(������   ;���   V�M��3���j �M�j/Q���  ��P����������Bd�H`jV�у���L���R���y���PW�������E�P�M�QWV�5����{@�C(�M�jV�������U�Rj���E�   �E�   �����������   ��U�R�Ћ���Qd�Bh�   V�Ћ{@�C(�M�jV�A�����V�M�������M��3���_^�   [�M�3��� ��]� _^3�[�M�3���� ��]� �M�^3�3�[��� ��]� ������������U���SV�uW�}�������u�����������H@�I�U�R�E�PW�ы]��E���UR�ΉE� ����EP�Ή]���������QH���  jW�Ѓ��MQ�ΉE���������Bd�W�у���t/����]�Bd�HXSW�у���t����Bd�HXSW�у������Bd�HW�у��؅�u����E������B@�@�M�Q�U�RS�ЋE���MQ�ΉE�>����U��EP�ΉU�-�����t����QH���  jS�Ѓ��E��E    �MQ��������M��  �UR�ΉE������E�P�M�Q�U�R�EP��� �  �MQ��������U�R�������E�P�������M�Q������_��^[��]������������SW��3�9_u萗  �G9_u`Vh�Oh�   h��j �aI  ����;�t5蓌  �������   ���   �҉F����F�F�^�^�^�w^�3��w���^������G(�_,�W �_�_8�G@�_D�_0_�   [� �V��W�~W��  ���N�    �;���_^� �������������U���$Vh'  �4  ����H�A�U�R�Ћ���Q�J�E�PV�ы���B�P<���M��҅�u����H�A�U�R�Ѓ��   ^��]�h�Oh  h��jH�=H  ������t����J  �4P�F    �F    �3�����Q�J�E�P�ы���B�Pj j��M�h�PQ�҃��E�P�M����  � V�M�QPj ��Rh�Y �P  ���M������  ����H�A�U�R�Ћ���Q�J�E�P�у���^��]���������U�조��P�B �� V��M$��=mric��   �NW3�;���   �ES�U$R�UP�ERP�}$�(����E�� �E�E��� W�E��F�P�WWR�E�P�U�RW�ŋ  �����]�3�3�;�t�P��X�U�P�U�P�U�P;V(u
;Nu�   3����}$���NQ�NQ��E�F�E�F �E�F$�V(�^,����B|�P����3��^8���F@�����FD�F0[;�tPPhI�����  ��_�   ^��]�  ����������U���T  SVW��� �}���  �����P�u���   ���$hxvpi�����]������Q���   ���$hyvpi�����]�����Q���   j hacpi���Ѓ��c  ��l������  �M����  �E�O�UR�UP�ERP�������_  �E��� �E��E��� j �E�G�P�j j R�E�P�U�Rj �#�  ��t+��O�P�w�V�H�N�P�V�H�N�P�u�V�!��G�X�E�@�����@    �     ���> ��  j h  ��  �E��]��j���\$���E��$h �  ��K  �E�P��T���Q��\���R���L  ���,  ���    ݅\���������������݅T�����Dz ����������Dz��j2�����  ����   �����E��U����E��U������ �E���� �j �E�G��@j j P�E�P�E�PR���  ��t"�;u�p�ыH�M̋H�MЋH�MԋH�����3��]�3�;O@u;W0u�   �3��W0�U�3ۅ��W4�U��ÉW8�UԉW<�O@�wD�Å�tj h%  �w�  ���u�]�E�P��T���Q��\���R����J  ����������K  ���  �G0;��  ����  ����P���   j haqpi�M��Ћ���O0�E䋂�   �Ph�  �҅���  �_0��������ˉE��������ˉu������؍M��]�>i  �E�j VSP�M��^i  �O0�^  �؉]����+  �
��$    �]�������   �Bh'  ���Ѕ���  �MSj(��  ��� �M�Q�E��U�R�U��E�P�E�M�QRVSP�ɤ �� 3ɉMЉMԉMظ    ��    �=�   r�;�t	P�M�������O(�W@�M��U��E�    ����   3��E��]�M�U�ۋ�������9��   3���$    ;�tq�M�ǃ�����;U�u[�M���Uċ�����Q�U�R�M̉E��w�����u)�Eč����Q��d���R�M̉�d���ǅh���    �����������M��H�E�G��|��}�@�E����H����E�@�E�;E�3����]�3�9u�>  �]��3��M�׃����U���9��   �M�������P�M�Q�M̉U����������� ��   ����ݕ����������ݕ����Qݕ����Vݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݝ����BD�U��@,R�Ћ������@3҃�;K�@��R�U��ʋ���̉�P�Q�P�Q�P�Q�P�@�Q�A������QW��������BD�U��@0������QVR�Ѓ�0G�������F��;u������}��]�������   �Bj j���ЍM�Q��;  �U�R��;  ���M�������E�P�E�    ��;  �u��������   �B(���ЉE���������M���e  ��  �E���K  �O0�w0j Q���f�  ���3  ��G(�ݕ<�����<���ݕD���RݕL���Pݕ$���Qݕ,����Mݝ4�����  ��؋G@��$���RPQ�M���ǒ  �W@�#؋G(RPQ�M貢  #��E�tT݅$����G@܅<����݅,���j ܅D����U�݅4���R܅L���P��PQ�M�����]������]����]�訒  #�3�;�tW��MWj"R�  ��tE�EP�j���V�d���W�	�  �MQ���  ���}�M����  ��l������  �   _^[��]� �UR谏  �}��EP袏  �E    ���M���  ��l�����  _^3�[��]� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������V����;  �<N��^�����������������;  �����������U��V����;  �Et	V�98  ����^]� ���������������U�조��Hd���   SV�uV�҃�P����Hd���   V�ҋu�]��P�E�P�����^[]��������������������������VW�q0�   ��    ������   ���V�҃�Oy�_^��������������������̋�3ɉ�H�H���̋A�������������V���X{  ���^�������������������V��V�G{  ���    ^������������̋�������������̋��������������V��V�{  ���    ^�������������U��E�]� ���̡��V�񋈈   ���   �҉��^��������������������̡��V�񋈈   ���   V�҃��    ^��������������̋�������������̋�������������̋�������������̋��     ��������V��V��  ���    ^������������̋�������������̋��������������V��V�Ǆ  ���    ^�������������U��E�]� ����U����M�]� �����������������̋�������������̋��������������U��E�]� ����3�9A����������V���X�  ���^�������������������V��V�W�  ���    ^������������̋�������������̋��������������U��E�	�@��]� �������������̃9 u�y ~�   �3��������������U��U���M��P]� �����������̋A�����������̋A������������̋��������������U��V�uV�#1  ���    ^]� ���������������������U����M���@    ]� ��������̋A�������������U�조��H�U����   �@h�N��j!P�у�]� ������������������U��V�u��MQ�E�{0  ���    ^]� �������������U���E� O��� ]� �����������U��E� �M3��1��]� �����������U�조��H�U����  hO��h5  P�у�]� �����������������̃9 u�y t�   Ãy ~�3�������̋��������������U���M��]� �����������������U��E]� ������U��E��U3�;
��]� ���������̋���������������U��E��t�M���Q�P�I�H]�3�]������������������������������U��U�E�V�2�0�
^]������������U��U�E�V�2�0�
^]�����������̋��     ������������������������U�조��UV�񋈄   �Aj RV�Ѓ���^]� ���������U��E��M;u�@;Au�   ]�3�]���������������U��E��u������A����]� ����R@V�qVQP�B�Ѓ�^]� ������������������������U��� �USV��W3��>�~�~�~�~ �~(����Hd���   �^h�  R�E�P�ы���}��}����   WP�A�U�R�Ћ�����   �
�E�P�ы�����   �PW�M�QV�ҡ�����   ��U�R�Ћ���Qd�E���   h�  P�M�Q�ҋ��W�}��}����   �JP�E�P�ы�����   ���D�M�Q�ҡ�����   W�U��ARS�Ћ�����   �
�E�P�ы���Bd�M���   jQ�U�R�Ћ��W�}��}����   �JP�E�P�ы�����   ��M�Q�ҡ�����   W�U�R�F P�A�Ћ�����   �
�E�P�у�@_��^[��]� ��������������������������������������������������������������������������������������������������������������������U��E��M;u�P;Qu�I;Hu�   ]�3�]�����������������������U��Uj j R�U����@P�ER�UPR�Lt  ]� ������������������������V���(2  �lO��^����������������2  �����������U��V���2  �Et	V�i.  ����^]� ���������������U��E�	�@��]� �������������̋A������������V��V��*  ���    �F    ^���������������������̋A�������������U��V�uW��9wu_�   ^]� ����H���  ShO��    h5  R�Ћ؃���tG��~C�G;�}�ƍ�    ���t��tQPS�t� ���G;�~��+���Q��j R��� ��W�*  ����w��t��u	[_3�^]� [_�   ^]� ������������������������������������������������������������������������U��E�U�RV�4���;�s)�UW��    ��t�:�9�z�y�z�y����;�r�_^]�������������������������������U��E]� ������U��E��U3�;
��]� ����������U���M��]� �����������������U��E�PV�q�p�Q�1��0�^]� ����������������U��E���]� ����������������U��Ej jP��z ��]������������U��EP�t(  ��]� �������������U����M�     ��P�I�H]� �������������������U��EV���u������F������^]� ����Q@�R�NQVP�҃���^]� �����������������U��VW�}���u3��F_������F������^]� ����H@�A�VRVW�Ћ���QH���  jW�Ѓ��F_��^]� �����������������������������������U��E�MW�x;yt3�_]�S3�V��~*�1� �N+��;u$�Y�;Xu�X;uB����;�|�^[�   _]�^[3�_]�����������������������3��A9A�����V��V��&  ���    �F    ^����������������������U��EV��P�    �F    �������^]� �������������U��S�]�V��;Fu^�[]� ����Q���   W�@h�N��j!P�ы�����t?��E�RQW��������~ ~��EP�U�&  ���    �>�_�N^�[]� _^2�[]� �������������������������������������U��QV��~ ~��M�Q�E��%  ���    �    �F    �F    ^��]��������������������U����EW��P�M��E�    �E�    �����}� uw�}� uwS3�9_~8V�W����t��F3��u��E��	�����0��u�G��    C;_|�^�E��O�G�E��W�G�E�P�M��U���$  ��[�   _��]� �}� ��M�Q��$  ��3�_��]� �����������������������������������������������������U��QV��FW�~;F}
��@���:@�E��E�� O��� �E��E�PW��������u_���^��]� ���@����t�M���Q�P�I�H��P�_^��]� �����������������������������������U��Ej jP�v ��]� ���������U��VW�}�7��t���E�u�6P�#  ����u��    _^]� ���������������U��E��t�M�     ��P�I�H]�3�]�������������U��QV��~ ~��M�Q�E��E#  ���    �    �F    �F    ^��]��������������������U��EVP�������> u�~ ~�   3Ʉ���^��]� 3�3Ʉ���^��]� �������������������3��A9A��   ���������������U��U��    ;�v�;�r�;AtP�$�����u]� �   ]� �������������U��SV��3�W9F��]�F;�t4�};�~-�E�EP�MQ��������u_^[]� �SWR�Ͼ�����~_^�[]� ������������������������U���W3��M�9y~5SV�A�4�����t�M��u��6Q��!  ����u�M�G�    ;y|�^[_��]����������������������U��Ej jP�s ��]� ���������U�조��H���  h�Mj{j�҃���t �M�     ��P�I�U�H�
�H]� �U�
3��H]� �������������������������������U���S�ك{ V�    �M�C    ������   ���   �sh�  j��E�    �Ѕ��   W�I ������   �E��M���   P�ҋ���u6����E�E��}�;C}U�@�������   �M��U��P�M�H�v����H@�I�U�R�E�PW�ы���BH���  jW�у��E��@�E��E�� O�� �U�RV�ˉE��������t!���@����t�U��M��H�U�P�����}����   �M���   h�  Gj��}���;�����_^[��]� �������������������������������������������������������������������������������������������̋�3ɉ�H�H����U��QV��~ ~��M�Q�E��%  ���    �    �F    �F    ^��]��������������������V���(f  �������   ���   �҉F����F�F3��F�F�F��^�������������������������V��读���F    ��V�  ���    �F    ^�����������������������U��QSV��3�W9^~�F�M�Q�E��A  ���^�^�^�^������   ���   �~W��V��be  ��_�^[��]�����������������������U��3�V��M�F�F�F�    ;�v	�I �;�r�;FtP���c�����^]� ����������������������U��Q�ES�VW�x��3��}9F��F;�t3;�~/�E��EP�M�Q���!�����u	_^[��]� �SWR�������~_^�[��]� ������������������������������U��S�]VWj ��~jS�8o 3����E�@    ����N���P��t�H�Q;t�H��P��u�_^3�[]� _^�   []� �����������������������������U��SVW�}j jW���n �ء���H���  h�Mj{j�҃���t�     ��H�W�P���3ɋ}�Y�O3ҋ��v�G    ��V������   F_^[]� ��������������������������������������������V��������F    ��V��  ���    �F    ^�����������������������U��3�V��M�F�F�F�    ;�v	�I �;�r�;FtP���#�����^]� ����������������������U���V��M�E�PQ��������E�U��0�P^��]� ����������������������U��QSV��3�W9^~�F�M�Q�E��  ���^�^�^�^������   ���   �~W��V��"b  ���E�t	V�  ��_��^[��]� �����������������������������������U��Q�ES�VW�x��3��}9F��F;�t6;�~2�E��EP�M�Q��������u_^��[��]� �SWR��������~_�^��[��]� ����������������������������������������U���VW�}�E�PW��蜶����u��U�E�R�E��M�P���	����E�M�_�0�H^��]� ���������������������������U��Q�ES�VW�x��3��}9F��F;�t*;�~&�E��EP�M�Q���!�����t�SWR�������~_��^[��]� �����������������������U��QSV�ً3W3�;�tc9~~�F�M�Q�E��  ���~�~�~�~������   ���   �~W��V�    �(`  V�    �  ��_^�    [��]É;_^[��]������������������������������������U��QSV�ً3W3�;�tc9~~�F�M�Q�E��k  ���~�~�~�~������   ���   �~W��V�    �_  V�    �l  ��_^�    [��]É;_^[��]������������������������������������U���VW�}�E�PW��茴����u��U�E�R�E��M�P��������E�M�_�0�H^��]� ���������������������������U��Q�ES�VW�x��3��}9F��F;�t*;�~&�E��EP�M�Q��������t�SWR� ������~_��^[��]� �����������������������V����  3��4P�F�F��^������̸�Y �����������U�조��H�QV�uV�ҡ���H�Qj j�h�PV�҃���^]� ��������������������������V��W�N�Ų���~W�h  ���    _��^�I  ���������U���VW�}�E�PW��������u��U�E�R�E��M�P���y����E�_��^��]� ����������������U��� ������   ���   SV��NW�ЋN�}jQ���?�  �E�UP�M�W3�Q��F�������B�}���   ��jh�  ���҉E���Ћ��S����� �с��   ��3��E
��3��S�]��с��   3��E��3��S�]�с��   ��3�3��S�]�M�NQ�M����������B���   j
h�  ���ҋ}��F9~u �FP�E�P�o�������t�M;Nu3���   �U�;��   �E�~�E9^�^�^9]�t2;�~.�EP�M�Q�N�]��z�����t�U��]�FRSP�b������^�M�U�R�N�E�P�M�Q�M�U�R�Z  ����}��]�+}�+]�Hd�U���   RGC�Ѓ��E    �t�E   �t�MV�[  ���    �s[  ���t9����Q�M���   j h�  �ЋM�V�6QPjR�URSW���[  ��u#�}� ~�E��MQ�E��  ��_^3�[��]� 3�9]�~�U��EP�U�  ��_^�   [��]� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������U��V��W�N�"����~W�e  �����    �  �Et	V�  ��_��^]� ����������������̡��V��H�QV�҃���^���������U�조��P�Rx]�����������������U�조��P�R@]�����������������U�조��P�RH]�����������������U�조��P�RL]����������������̋�������������̡�����   �BHQ�Ѓ������������̡�����   �BTQ�Ѓ�������������U�조��P�E���   ��VWP�EP�E�P�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ������������U��E��u����MP�EPQ��  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h�Pj;h��j��  ����t
W����  �3��F��u_^]� �~ t3�9_��^]� ����H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ����H<�Q��3Ʌ����^��������������̃y t�   ËA��uË���R<P��JP�у��������U����u����H�]� ����J<�URP�A�Ѓ�]� ���������������U�졠���u����H�]Ë���J<�URP�A�Ѓ�]�U�졠���$V��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�SP�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���[t.����B�u�HV�ы���B�P�M�Q�҃���^��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^��]���������������U�졠���$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]����������������U�졠���$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]��U�졠���$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hQP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]����U�조��H<�A]����������������̡���H<�Q�����V��~ u>���t����Q<P�B�Ѓ��    W�~��t�����  W�4	  ���F    _^��������U���V�E�P���N�  ��P�������M����  ��^��]��̃=�� uK�����t����Q<P�B�Ѓ����    �����tV���p�  V�  �����    ^������������U���H����H�AS�U�V3�R�]��Ћ���Q�JSj��E�hQP�ы���B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]�� �M�Q�U�R�M��� ���&  W�}�}���   ������   �U��ATR�Ћ�������   ����Q�J�E�P���ы���B���   ���M�Qj�U�R���Ћ���Q�J���E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Bx��W�M����E���t�E� ��t����Q�J�E�P����у���t����B�P�M�Q����҃��}� u"�E�P�M�Q�M���  ��������E�_^[��]ËU��U�_�E�^[��]��U���DSV�u3ۉ]�;�u_����H�A�U�R�Ћ���Q�JSj��E�hQP�ы���B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]����  �M�Q�U�R�M��1  ���p  W�}��I �E����   ������   �U��ATR�Ћ�������   ����Q�J�E�P���ы���B���   ���M�Qj�U�R���Ћ���Q�J���E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Bx��W�M����E��t�E ��t����Q�J�E�P����у���t����B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*������   P�BH�Ћ���Q���ȋBxW�Ѕ�t"�M�Q�U�R�M����  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��3�  �EP�M�Q�M�u��u�}�  ����   �u���E���tA��t<��uZ������   �M�PHQ�ҋ���Q���ȋBxV�Ѕ�u-�   ^��]Ë�����   �E�JTP��VP�[�������uӍUR�E�P�M����  ��u�3�^��]����������V��~ u>���t����Q<P�B�Ѓ��    W�~��t���z�  W�  ���F    _^��������U��V���U�  �Et	V�  ����^]� ���������������U�조��P�E�RxP�����@]� ���U��E���� ]��U��V�u���t����QP��Ѓ��    ^]���������̡���H��@  hﾭ���Y����������U��E��t����QP��@  �Ѓ�]����������������U�조��H���  ]��������������U�조��H��  ]�������������̡���H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW膪 ������u_^]Ã} tWj V蜠 ��_������F���   ^]���U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�
� ������u_^]�Wj V�&� ��_������F���   ^]�������������U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW芩 ������u_^]�Wj V覟 ��_������F���   ^]�������������U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�
� ������u_^]�Wj V�&� ��_������F���   ^]�������������U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW芨 ������u_^]�Wj V覞 ��_������F���   ^]�������������U��M��t-�=�� t�y���A�uP��� ��]á���P�Q�Ѓ�]��������U��M��t-�=�� t�y���A�uP耨 ��]á���P�Q�Ѓ�]��������U�조��H�U�R�Ѓ�]���������U�조��H�U�R�Ѓ�]���������U�����E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�F� ������u_^]�Wj V�b� ��_������F���   ^]���������U�����E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]Ã�s�   VW�xW蝦 ������u_^]Ã} tWj V賜 ��_������F���   ^]����������U��E��u�   �����t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�� ������u_^]�Wj V�3� ��_������F���   ^]����������U��E��u�   �����t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW脥 ������u_^]�Wj V蠛 ��_������F���   ^]�������U�조��H�U�R�Ѓ�]���������U�조��H�U�R�Ѓ�]���������U�조��H�U�R�Ѓ�]���������U�조��H�U�R�Ѓ�]��������̋��  Q��������� Q���������̅�t��j�����̡���P��  �ࡰ��P��(  ��U�조��P��   ��V�E�P�ҋuP����  �M����  ��^��]� ��������̡���P��$  ��U�조��H��  ]��������������U�조��H���  ]�������������̡���H��  ��U�조��H���  ]��������������U�조��H��x  ]��������������U�조��H��|  ]�������������̡���H��d  ��U�조��H��p  ]��������������U�조��H��t  ]��������������U���EV��� Qt	V���������^]� ��������������U��E#E]������U��E#E]�����̋A������������̸   � ��������� ������������̃��� ����������� �������������U�조��H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ����Q0�F�M���   PQW�ҋF��^_]� U�조��H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U�조��H���  ]��������������U�조��H���  ]��������������U�조��P�EP�EP�EP�EPQ���   �у�]� �����U�조��E�P�EP�E���\$�E�$PQ���   �у�]� �������������U�조��P�EP�EP�EPQ���   �у�]� ��������̡���P���   Q�Ѓ�������������U�조��P�EP�EP�EPQ���   �у�]� ���������U�조��P�EP�EPQ���   �у�]� �������������U�조��H�U�ApR�Ѓ�]� �����U�조��P�EP�EPQ���  �у�]� �������������U�조��P�EP�EPQ���  �у�]� �������������U�조��P�EP�EPQ���  �у�]� �������������U�조��P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P贔 ��R���E�P���ҡ���P�B<�M��Ћ}��t0j �M�QW�q�������u����B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4���p} �E��� �E�Ї �E�0� �E��� �E��� �E��� �E�� ǅx���`� ǅ|���p� �E��� �E�@� �E�P� �E��� �E�P� �E�`� �E��� �E� � �E� � �E��� �E�p� 踋  ������B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u����H�A�UR�Ѓ�^3�[��]Ë���Q�B<W�M3��Ѕ��N  ���  �E�����   �MQ�M���  ����B�P�M�Q�ҡ���H�AWj��U�h$QR�Ѓ��M�Q�M��{�  �u�Wj��U�R�E�P��\���Q�_?�^�  ��P��x���R�n�  ��P�E�P�a�  ��P����  �E���t�E� �� t�M������  ��t��x��������  ��t��\�������s�  ��t�M̃���c�  ��t����Q�J�E�P����у���t�M��9�  �}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R��  ����E$�M�UVP�Ej QRP�������������Q�J�EP�у���_^[��]���������U��E�M�UP�EQ�Mj RPQ������]��������������V���(�  ���^���V��V�'�  ���    ^������������̋�������������̋�������������̋�`<����������̋�`L����������̋�`����������̋�` ����������̋�`0����������̋�`P����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`����������̋�`����������̋�`,�����������U��E��E	]�̋�3ɉ�H�H�H�H�H�H��������U�조��P�B4VW�}j��h�  ���ЋMWQ������_^]� ��������������U��V���PXW�ҋ}P����  ���Et�_�   ^]� �M�UPWQR������_^]� �����������U��S�]VW��j ���|�  �8�  �}uI�~ uC����P���   j h�  ���Ѕ�u����QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ������_^[]� ��������U��EP�A    �-�  ��]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �y  ����   �M3�V芲  �8�  u4��v  P�w�  ����P�M�B4��jh�  ��_^�C�[��]� �MV�E�  �8�  u�E�M��RPQ����_^�   [��]� �MV��  �8�  t�MV��  �8��  ����P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P�����3��؃��u�;�t����QH���  VS�Ѓ��E��M�;O�b  9w�Y  ����B�M���   Vh�  �҅�u!����P�M���   Vh�  �Ѕ��  ����Q�M�B4Vh�  ��;�t
V���������E��G������   ���   �Ћ]�E�;���   ;���   S�W}  �M���jQ�ˉu��uĉuȉủuЉu؉u��b  �U�E��ˉu��u�u�U�E��]��E�   ��q  ��tHtHt�u���E�   ��E�   ��E�   ��  �M�;�t�2v  ��BX�M�Q����P�߅  �M܃�;�t�0v  �M��X�  �M��P�  �M��R����]�U�E�MRSPQ���Q���_^[��]� ������   ���   �E�P�у�_^�   [��]� ���������������h��Ph:� �@�  ���������������U��Vh��jh:� ����  ����t�@��t�MQV�Ѓ�^]� ���^]� ����U��Vh��jh:� �����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh��jh:� ����  ����t&�@��t�M�UQ�MR�UQ�MRQV�Ѓ�^]� 3�^]� �����U��Vh��jh:� ���I�  ����t"�@��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��h��j h:� ���  ����t
�@ ��t]��3�]��������U��h��j$h:� ���  ����t
�@$��t]��3�]��������U��Vh��j(h:� ����  ����t"�@(��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh��j,h:� ���I�  ����t�@,��t�MQV�Ѓ�^]� 3�^]� �����U��M�E;�|	�E;���]���������U���E�E������{���E������z��]���]���������U�조��P�E���   ��P�EP�E�P�ҋM���P�Q�P�Q�P�Q�P�@�Q�A����]� �U�조��E�P�E�R,���$P��]� ���������������U�조��P�RH]����������������̡�����   �B��U�조����   �RH]��������������U�조��P@�EP�EPQ�J(�у�]� ����P@�B,Q�Ѓ���������������̡���P@�B,Q�Ѓ���������������̡�����   �Bx��U�조����   �R|]�������������̡�����   �B(��U�조��PH�EP�EPQ���   �у�]� �������������U�조��PH�EP�EPQ���   �у�]� �������������U�조��PH�EPQ���   �у�]� �U�조��PH�EPQ���   �у�]� �U�조��PH�EPQ���   �у�]� ̡���PH���   j h�  Q�Ѓ�����̡���PH���   j h(  Q�Ѓ�����̡���PH���   h(  Q�Ѓ�������̡���PH���   j h�  Q�Ѓ������U�조��Pl�E�I�RP�EP�EP�EPQ�҃�]� �����U�조��Pl�E�I�RPQ�҃�]� �U�조��P\�EPQ�J,�у�]� ���̋���Ѓ������̋��%��������̋A�������������U���M����%���]� ���������U���M�����Ѓ�]� ��������̃y ~�� ��%���Ã������������U�조��E�PH�B���$Q�Ѓ�]� ���������������U�조��PH�EPQ���   �у�]� �U�조��PH�EPQ���  �у�]� �U�조��PH�EPQ���  �у�]� �U�조��PH�EP�EPQ��  �у�]� �������������U�조��PH�EP�EPQ��  �у�]� ������������̡���PH���  Q�Ѓ�������������U�조��PH�EPQ���  �у�]� ̡���PH���   j Q�Ѓ�����������U�조��PH�EPj Q���   �у�]� ��������������̡���PH���   jQ�Ѓ�����������U�조��PH�EPjQ���   �у�]� ��������������̡���PH���   jQ�Ѓ����������U�조��PH�EPjQ���   �у�]� ���������������U�조��PH�EP�EPQ���   �у�]� �������������U�조��PH�EP�EPQ���   �у�]� ������������̡���PH���   Q�Ѓ�������������U�조��PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���0�  ������t�E����QH���   PVW�у���_^]� �����U��EVW���MPQ�<�  ������t�M����BH���   QVW�҃���_^]� ̡���PH���   Q�Ѓ������������̡���PH���   Q�Ѓ�������������U�조��PH�EPQ���   �у�]� �U�조��PH�EPQ���   �у�]� �U�조��PH�EP�EPQ��8  �у�]� �������������U�조��PH�EP�EPQ��   �у�]� ������������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ������������̡���PH��  Q�Ѓ������������̡���PH��  Q�Ѓ�������������U�조��PH�EP�EPQ��  �у�]� �������������U�조��PH�EP�EP�EPQ��   �у�]� ���������U�조��PH�EP�EP�EP�EPQ��|  �у�]� �����U�조��PH�EPQ��  �у�]� ̡���PH��T  Q�Ѓ�������������U�조��PH�EP�EPQ��  �у�]� �������������U�조��PH�EPQ��8  �у�]� �U�조��PH�EPQ��<  �у�]� �U�조��PH�EP�EP�EPQ��@  �у�]� ���������U�조��PH�EPQ���  �у�]� ̡���PH��L  Q��Y��������������U�조��PH�EPQ��H  �у�]� ̡��V��H@�Q,WV�ҋ���Q��j �ȋ��   h�  �Ћ���QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡���P@�B,Q�Ћ���Q��j �ȋ��   h�  �������U�조��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�조��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�조��PH�EP�EP�EPQ��   �у�]� ��������̡���HH��  ��U�조��HH��  ]��������������U�조��E�PH��$  ���$Q�Ѓ�]� �����������̡���PH��(  Q�Ѓ�������������U�조��PH�EP�EPQ��,  �у�]� �������������U�조��E�PH�EP�E���$PQ��0  �у�]� ���̡���PH���  Q�Ѓ������������̡���PH��4  Q�Ѓ������������̋��     �������̡���PH���|  jP�у���������U�조��UV��HH��x  R��3Ƀ������^��]� ��̡���PH���|  j P�у��������̡���PH��P  Q�Ѓ������������̡���PH��T  Q�Ѓ������������̡���PH��X  Q�Ѓ�������������U�조��PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡���PH��`  Q�Ѓ�������������U�조��PH�EPQ��d  �у�]� �U�조��E�PH��h  ���$Q�Ѓ�]� ������������U�조��E�PH��t  ���$Q�Ѓ�]� ������������U�조��E�PH��l  ���$Q�Ѓ�]� ������������U�조��PH�EPQ��p  �у�]� �U�조��PH�EP�EP�EP�EPQ���  �у�]� �����U�조��PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U�조��E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E����HH�E���   R�U���$P�ERP�у�]����������������U���E�M�(Q�l} �M;�|�M;�~��]�����������U�조��PH�E���   Q�MPQ�҃�]� ������������̡���PH���   Q��Y�������������̡���PH���   Q�Ѓ������������̡���PH���   Q��Y��������������U�조��PH�EP�EPQ���   �у�]� �������������U�조��PH�EP�EP�EP�EP�EPQ���  �у�]� ̡���PH��t  Q��Y�������������̋�� <Q�@    ��<Q����Pl�A�JP��Y��������U�조�V��Hl�V�AR�ЋE����u
�   ^]� ����Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË���QlP�B�Ѓ�������U�조��Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E����HH�ER�U���$P���  R�Ѓ�]����U�조��HH���  ]��������������U�조��HH���  ]��������������U��U0�E(����HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U�조��HH���  ]��������������U�조��E�PH�EP���$Q���  �у�]� ��������U���V�����  �E����   �} ��   ����HH��p  SWj h�  V�ҋء���HH���   h�  V�]��ҋ������}����   �M3��u���  ����   �]�E�P�M�Q�MWV�z�  ��t\�u�;u�T������u�E����ҋL�;L�t-����Bl�S�@����QR�ЋD������t	�M�P�c�  F;u�~��}�u�MF�u��+�  ;��w����E�_[^��]� 3�^��]� ��������������U������SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u����HH���  �'��u����HH���  ���uš���HH���  S�ҋȃ��E��t�W���  ����HH���   h�  S3��҃����  ���_�u����    ����Hl�U�B�IWP�ы�������   ����F�J\�UP�A,R�Ѓ���t�K�Q�M��  ����F�J\�UP�A,R�Ѓ���t�K�Q�M���  �E��;Pt&�F����Q\�J,P�EP�у���t	�MS��  ����v�B\�M�P,VQ�҃���t�M�CP��  ����QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U�조��HH���   ]�������������̡���PH���   Q��Y��������������U�조��HH���  ]��������������U�조���P���   V�uW�}���$V�����E������At���E������z����؋���Q�B,���$V����_^]����������������U���0���U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١���]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U�조��HH�]��U�조��H@�AV�u�R�Ѓ��    ^]�������������̡���HH�h�  �҃�������������U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��HH�Vh  �ҋ�������   �EPh�  �`�  ����t]����QHj P���   V�ЋMQh(  �6�  ����t3����JH���   j PV�ҡ�����   �B��j j���Ћ�^]á���H@�QV�҃�3�^]�������U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��HH�Vh�  �ҋ�����u^]á���HH�U�E��  RPV�у���u����B@�HV�у�3���^]�������U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��HH�I]�����������������U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��PH�EPQ���  �у�]� �U�조��PH�EPQ���  �у�]� ̡���PH���  Q�Ѓ�������������U�조��HH���  ]��������������U�조��E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡���PH���  Q�Ѓ�������������U�조��PH�EP�EPQ���  �у�]� ������������̡���PH��  Q�Ѓ�������������U�조��PH�EP�EP�EPQ���  �у�]� ��������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ�������������U�조��PH�EPQ��  �у�]� �U�조��PH�EPQ��  �у�]� ̋������������������������������̡���HH���  ��U�조��HH���  ]��������������U�조��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U�조��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡���PH��,  Q�Ѓ�������������U�조��PH�EPQ��X  �у�]� ̡���PH��\  Q�Ѓ�������������U�조��HH��0  ]��������������U�조���W���HH���   j h�  W�҃��} u�   _��]� Vh�  �߆  ��������   ����HH���   j VW�҃��M���  ����P�E�R0Ph�  �M����E����P�B,���$h�  �M��Ћ���Q@�J(j �E�PV�у��M���  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7����U�HH���   RW�Ѓ���u����QH���   jW�Ѓ���t�   �����   ����QH���   W�Ѓ��} u(����E�QH�M���  P�ESQ�MPQW�҃��B�u��t;����U�HH�ER�USP���  VRW�Ћ�����   �B(�����Ћ���uŃ; u����QH���   W�Ѓ���t3���   �W��u1����QH���   �Ћ���E�QH���   PW�у�_^[]� ����BH���   �у��} u0����M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ����QH�h  �Ћ؃���u_^[]� ������   �u�Bx���Ћ�����   P�B|���Ѕ�tU����E�QH�MP�Ej Q���  VPW�у���t������   �ȋBHS�Ћ�����   �B(���Ћ���u�_^��[]� ��������������U��EV���u����HH���  �'��u����HH���  ���u����HH���  V�҃���u3�^]� P�EP���.���^]� ���������U���D����HH���   S�]VWh�  S�ҋ���HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��>
  ������   �B���Ћ��=�  �  �QH���   Wh:  S�Ћ���QH�E����   h�  S�Ћ���QHW�����   h�  S�uԉ}��Ћ���QH�E苂  S�Ћ���QH�EЋ��  S�Ѓ�(�E��E�HQ��~~�M���M�I �MЅ�tMj�W��  ���t@�@�Ẽ|� �4�~����%�������;�u/�����  ;E�~�E؋���  E���E�;Pu�E���E��E�G;}�|��}� ��   �u�j S���ׁ  ����  ���ȅ  ��ti���m  �}�;�u^����H���  �4�hLQ��h�  V�҃��E���b  �M��E��y�  ��t�}� t��tVP�E�P� f ����}܋���Q���  �4�hLQ��h�  V�Ѓ��E����  �M�3�;�t;�tVQP�e ���E�;�~-����QhLQ��h�  P���   �Ѓ��E�;���  ����E��QH��  j�PS�у�����  �u�;�tjS��襀  ���{  ��趄  �E���}����BH���   Wh�  S�у�3��E�}�9}��]  �}���}����$    �MЅ��J  �U�j�R��  ����6  �M̍@�|� ���]�~����%�������9E���  ���m�  �E�3�3ɉE܉M�9C��   ��$    �����������ti�]������������M�ҋ9�<��}�҉T��y�]��|��]��z�|��y�]��|��]��z�|��I�}��]��L��M��}ȃ��T����M�A�M�;K�v����E؅��0  �+U�j��PR�M����  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t4�U�M��@���P�Q�P�Q�P�Q�P�Q�@�A�M��Eȍ@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A;]�}_�UȋE�9�uT�ȋL�����������w0�$�d� �U���4���M���t���U���t��	�M���t��M���;]�|��E܃�F�M�;]������U�;U��  �U�R�y����E�P�p����M�Q�g�����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q�P �Q�P$�Q�P(�I�H,��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@���E��}�;E�������U�R�\����E�P�S������  ���   �B����=  ��  ����QH���   j h(  S�Ћ���QH�����   h(  S�ЋЃ�3��U؅�~"��ǅ�t�|� t�4N��tN�@;�|�u��u܋���Q���  �4v�hLQ��hK  V�Ѓ��E�����   �M��t��tVQP��_ ���u؋���Q���  �hLQ��hP  V�Ѓ��E���tP��t��tVWP�_ ���M����+���RH��PQ�E���   S�Ѓ���u�M�Q�����U�R�	�����_^3�[��]á���HH���   j h�  S�҉E�����HH���   j h(  S��3�3���3��E��}ĉ]�9]��:  �U��څ��  �E�    ����   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T�Y�Z�Y �Z�Y$�Z�Y(�R�]��Q,�U�@����0��;�|��}ă|� �t   �U��M�ύI�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�Tv�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}�C�]�;]�������M�3�3�;�~�U���$    �t���   @;�|��U�R�G������E�P�;�����_^�   [��]û� ŵ е ۵ �����������̋�� 4Q��������U��U��t�M��t�E��tPRQ� ] ��]������������U��U��t�M��t�E��tPRQ��\ ��]�����������̋�� HQ��������U��E� �M+]� ���������������U��V��V�<Q����Hl�AR�Ѓ��Et	V脽������^]� ����������U����M�3ɉH�H]� ����������U�조��Hd�IP]�����������������U��E�8 t����QdP�BT�Ѓ�]��U�조��Ph�EP�EP�EP�EPQ�
�у�]� ���������U�조��Ph�EP�EP�EP�EPQ���   �у�]� �����U�조��Ph�EP�EP�EPQ�J�у�]� ������������U�조��Ph�EP�EP�EP�EP�EPQ�J �у�]� ����U�조��Ph�EP�EP�EP�EPQ���   �у�]� �����U�조��Ph�EPQ���   �у�]� ̡���Hh�QX�����U��E�8 t����QhP�B\�Ѓ�]��U�조��Ph�E P�EP�EP�EP�EP�EP�EPQ�J`�у� ]� ������������U�조��Ph�E P�EP�EP�EP�EP�EP�EPQ�Jd�у� ]� ������������U�조��Ph�EP�EPQ�Jh�у�]� U�조��Ph�EP�EPQ�Jl�у�]� U�조��Ph�EP�EPQ�Jp�у�]� U�조��Ph�EP�EP�EPQ�Jt�у�]� ������������U�조��Hh���   ]��������������U�조��Ph�EPQ�Jx�у�]� ����U�조��Ph�E P�EP�EP�EP�EP�EP�EPQ���   �у� ]� ���������U�조��Ph�E P�EP�EP�EP�EP�EP�EPQ���   �у� ]� ���������U�조��Ph�E P�EP�EP�EP�EP�EP�EPQ���   �у� ]� ���������U�조��Ph�EP�EP�EPQ�J|�у�]� ������������U�조��E�Ph�E P���\$�E�\$�E�$Q���   �у� ]� ����������U�조��Ph�EP�EP�EP�EP�EPQ���   �у�]� �U�조��Ph�EP�EP�EP�EPQ���   �у�]� �����U�조��Hh���   ]��������������U����EV�uW���M�Q�M��    �F    �E��E�    �E�    ��  j V�U�R����  �M��z  _��^��]� ������U�조��E�Ph�EP���$Q���   �у�]� ��������U�조��E�Ph�EP���$Q���   �у�]� ��������U�조��Ph�EP�EPQ���   �у�]� �������������U�조��Ph�EP�EPQ���   �у�]� �������������U�조��E�Ph�E(���   ��P�E$P�E���\$�E�$P�EPQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A��(����]�$ �����U�조��E�Ph�E$���   ��P�E���\$�E�$P�EPQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A��$����]�  ���������U�조��P�Rp]�����������������U�조����   �R@]��������������U�조����   �RD]�������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t������   P�B@��]� �E��t������   P�BD��]� ������   R�PD��]� �����U�조��P@�Rd]�����������������U�조��P@�Rh]�����������������U�조��P@�Rl]�����������������U�조��P@�Rp]�����������������U�조����   ���   ]�����������U�조����   ���   ]����������̡���P@�Bt����̡���P@�Bx�����U�조��P@�R|]����������������̡���P@���   �ࡰ����   �Bt��U�조��P@���   ]�������������̡���P@���   ��U�조��P@���   ]��������������U�조��P@���   ]��������������U�조��P@���   ]��������������U�조��P@���   ]��������������U�조��P@���   ]��������������U�조��P@���   ]��������������U�조�V��H@�QV�ҋM����t��#�������Q@P�BV�Ѓ�^]� �̡���PH���   Q�Ѓ�������������U�조��P@�EPQ�JL�у�]� ���̡���P@�BHQ�Ѓ����������������U�조��P@�EP�EP�EPQ�J�у�]� ������������U�조��P@�EPQ�J�у�]� ����U�조��P@�EP�EPQ�J�у�]� U�조��P@�EPQ�J �у�]� ����U�조����   �R]��������������U�조����   �R]��������������U�조����   �R ]��������������U�조����   ���   ]�����������U�조����   ��D  ]�����������U�조��E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U�조����   ���   ]����������̡�����   �B$�ࡰ��H@�Q0�����U�조��H@�A4j�URj �Ѓ�]����U�조��H@�A4j�URh   @�Ѓ�]�U�조��H@�U�E�I4RPj �у�]�̡���H|�������U��V�u���t����Q|P�B�Ѓ��    ^]��������̡���H|�Q �����U��V�u���t����Q|P�B(�Ѓ��    ^]��������̡���H@�Q0�����U��V�u���t����Q@P�B�Ѓ��    ^]���������U�조��H@���   ]��������������U��V�u���t����Q@P�B�Ѓ��    ^]��������̡���PH���   Q�Ѓ�������������U�조��PH�EPQ��d  �у�]� �U�조��H �IH]�����������������U��}qF uHV�u��t?������   �BDW�}W���Ћ���Q@�B,W�Ћ���Q�M�Rp��VQ����_^]����������̡���P@�BT�����U�조��P@�RX]�����������������U�조��P@�R\]����������������̡���P@�B`�����U�조��H��T  ]��������������U�조��H@�U�A,SVWR�Ћ���Q@�J,���EP�ы���Z��h��hE  �΋���e  Ph��hE  ����e  P��T  �Ѓ�_^[]����U����M�]� ��U��U���M��P]� ������������U����M�]� ��U����M�]� ��h��Ph� 蠽  ���������������h��jh� ��  ����uË@����U��V�u�> t/h��jh� �S�  ����t��U�M�@R�Ѓ��    ^]���U��Vh��jh� ����  ����t�@��t�M�UQR����^]� 3�^]� ���U��Vh��jh� ���ټ  ����t�@��t�M�UQR����^]� 3�^]� ���U��Vh��jh� ��虼  ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������Vh��jh� ���L�  ����t�@��t��^��^��������U��Vh��j h� ����  ����t�@ ��t�MQ����^]� ��������������U��Vh��j$h� ���ٻ  ����t�@$��t�M�UQR����^]� 3�^]� ���U��Vh��j(h� ��虻  ����t�@(��t�M�UQR����^]� 3�^]� ���U��Vh��j,h� ���Y�  ����t�@,��t�M�UQR����^]� 3�^]� ���U��Vh��j0h� ����  ����t�@0��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��j4h� ���ɺ  ����t �@4��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��j8h� ���y�  ����t%�@8��t�M�E�UQ�M���$RQ����^]� 3�^]� ������U��Vh��j@h� ���)�  ����t�@@��t�M�UQR����^]� 3�^]� ���U��Vh��jDh� ����  ����t�@D��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jHh� ��虹  ����t �@H��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��jLh� ���I�  ����t�@L��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jPh� �����  ����t�@P��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jTh� ��詸  ����t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��jXh� ���Y�  ����t �@X��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��jdh� ���	�  ����t%�@d��t�E�M�U���$Q�MRQ����^]� 3�^]� ������U��Vh��jhh� ��蹷  ����t �@h��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��jlh� ���i�  ����t$�@l��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh��jph� ����  ����t �@p��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��jth� ���ɶ  ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vh��jxh� ��艶  ����t �@x��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh��j|h� ���9�  ����t�@|��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��h�   h� ����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h� ��薵  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h� ���F�  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h� �����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h� ��覴  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h� ���V�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ��足  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h� ���f�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���Ʋ  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���v�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���&�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���ֱ  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h� ��膱  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��j\h� ���9�  ����t�@\��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��j`h� ����  ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vh��j<h� ��詰  ����t$�@<��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh��h�   h� ���V�  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   h� ����  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   h� ���֯  ����t'���   ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh��h�   h� ��膯  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���6�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h� ��薮  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���F�  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h� �����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ��覭  ����t,���   ��t"�E�M�U���$Q�MR�UQR����^]� 3�^]� ������������U��Vh��h�   h� ���F�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� �����  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h� ��覬  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ���V�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   h� ����  ����tG���   ��t=�E(�MP���ĉ�M�H�M�H�M�H�M �H�M$�H�E�MPQ����^]�$ 3�^]�$ �U��Vh��h�   h� ��薫  ����tN���   ��tD�E0�E(�MP�� ���\$��M�H�M�H�M�H�M �H�M$�H�E�MPQ����^]�, 3�^]�, ����������U��Vh��h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h   h� ���ƪ  ����t��   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h  h� ���v�  ����t#��  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h  h� ���&�  ����t��  ��t�M�UQR����^]� 3�^]� �������������U��Vh��h  h� ���֩  ����t��  ��t�M�UQR����^]� 3�^]� �������������U��Vh��h  h� ��膩  ����t'��  ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh��h  h� ���6�  ����t#��  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h  h� ����  ����t'��  ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh��h  h� ��薨  ����t��  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h   h� ���F�  ����t��   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h$  h� �����  ����t#��$  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h(  h� ��覧  ����t#��(  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h,  h� ���V�  ����t3��,  ��t)�M$�U Q�MR�UQ�MR�UQ�MR�UQR����^]�  3�^]�  �����U��Vh��h0  h� �����  ����t��0  ��t�MQ����^]� ��������U��Vh��h4  h� ��趦  ����t��4  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h8  h� ���f�  ����t��8  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h<  h� ����  ����t#��<  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h@  h� ���ƥ  ����t#��@  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��hD  h� ���v�  ����t��D  ��t�M�UQ�MRQ����^]� U��Vh��hH  h� ���6�  ����t��H  ��t�M�UQ�MRQ����^]� U���V��FT��u
���^��]� �V$�MjRP�E�M�P�M��E��Q膭  ��t�+FT^����]� �����U���V��FX��u
���^��]� �V(�MjRP�E�M�P�M��E��Q�6�  ��t�+FX^����]� �����U���V��F\��u
���^��]� �V,�MjRP�E�M�P�M��E��Q��  ��t�+F\^����]� �����U���V��FL��u
���^��]� �V4�MjRP�E�M�P�M��E��Q�E�����菬  ��t�+FL^����]� ��������������U���V��F<��u
���^��]� �V$�MjRP�E�M�P�M��E��Q�6�  ��t�+F<^����]� �����U���V��F@��u
���^��]� �V(�MjRP�E�M�P�M��E��Q��  ��t�+F@^����]� �����U���V��FD��u
���^��]� �V,�MjRP�E�M�P�M��E��Q薫  ��t�+FD^����]� �����U���V��FP��u
���^��]� �V �MjRP�E�M�P�M��E��Q�F�  ��t�+FP^����]� �����U���V��FH��u
���^��]� �V0�MjRP�E�M�P�M��E��Q�E�������  ��t�+FH^����]� ��������������U���V��F8��u
���^��]� �V �MjRP�E�M�P�M��E��Q薪  ��t�+F8^����]� ����̋�� �Q��������U��E� �M+]� ��������������̋�� �Q��������U��E�@�M+A]� ������������̋�� �Q��������U��E� �M+]� ���������������U��EE]�������������X�����U���E���X�    ]� �����������U����M�    �H]� �����������U��UV���    �F    ������   �A(RV�Ѓ���^]� ��������������U��UV���    �F    ������   �A,RV�Ѓ���^]� �������������̡�����   �B8Q�Ѓ������������̡�����   �B<Q�Ѓ������������̡�����   �BLQ�Ѓ������������̡�����   �BPQ�Ѓ�������������U�조����   �R]��������������U�조����   �R<]�������������̡�����   �BP�ࡰ��HL���   ��U�조��H@�AV�u�R�Ѓ��    ^]�������������̡���HL�������U�조��H@�AV�u�R�Ѓ��    ^]�������������̡���PL���   Q�Ѓ�������������U�조��PL�EP�EPQ���   �у�]� �������������U�조�V��HL���   V�҃���u����U�HL���   j RV�Ѓ�^]� ������   �ȋBP�Ћ�����   �MP�BH��^]� �����̡���PL��(  Q�Ѓ�������������U�조��PL�EP�EPQ��,  �у�]� ������������̡���HL�Q�����U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��PL�E�R��VPQ�M�Q�ҋu��P���%D  �M��=D  ��^��]� ����U�조��PL�EPQ���   �у�]� �U�조��PL�EP�EPQ�J�у�]� ����PL�BQ�Ѓ���������������̡���PL�BQ�Ѓ���������������̡���PL�BQ�Ѓ����������������U�조��PL�EP�EP�EPQ�J �у�]� ������������U�조��PL�EPQ��4  �у�]� �U�조��PL�EP�EP�EPQ�J$�у�]� ������������U�조��PL�EP�EP�EP�EPQ�J(�у�]� �������̡���PL�B,Q�Ѓ���������������̡���PL�B0Q�Ѓ����������������U�조��PL�EP�EPQ��  �у�]� ������������̡���PL���   Q�Ѓ�������������U�조��PL�E��  ��VPQ�M�Q�ҋu��P���B  �M��B  ��^��]� ̡���PL�B4Q�Ѓ���������������̡���PL�B8j Q�Ѓ��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL��l  ]��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL���   ]��������������U�조��PL�EPQ�J<�у�]� ���̡���PL�BQ��Y�U�조��PL�EP�EPQ�J@�у�]� U�조��PL�Ej PQ�JD�у�]� ��U�조��PL�Ej PQ�JH�у�]� ��U�조��PL�EjPQ�JD�у�]� ��U�조��PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}���X  W�M�Q�U�R���������M�����J  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �X  j�M�Q�U�R�������M��J  ������   ��U�R�Ѓ�^��]�����������U���$����UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��W  j�E�P�M�Q�������M��I  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��W  j�E�P�M�Q�������M��I  ������   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��V  W�M�Q�U�R���������M����H  ��t+�u����[  ������   ��U�R�Ѓ�_��^[��]� ������   �JL�E�P�ыu��P���E\  ������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���U  W�M�Q�U�R����������M�����G  ��t+�u���[  ������   ��U�R�Ѓ�_��^[��]� ������   �JL�E�P�ыu��P���[  ������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��4U  W�M�Q�U�R���������M����'G  _^��[t������   ��U�R�������]Ë�����   �J<�E�P���]�������   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��T  W�M�Q�U�R���d������M����wF  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}���S  W�M�Q�U�R���������M�����E  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� �����̡���PL���   Q��Y��������������U�조��PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U�조��PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��DR  W�M�Q�U�R���$������M����7D  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��tQ  W�M�Q�U�R���T������M����gC  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��P  W�M�Q�U�R���������M����B  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���O  W�M�Q�U�R���������M�����A  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �O  j�M�Q�UR�������M�A  ������   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��N  j�U�R�E�P�������M��@  ������   �
�E�P�у�^��]� ��������U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��*N  j�E�P�M�Q���)����M��!@  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��M  j�E�P�M�Q�������M��?  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��*M  j�E�P�M�Q���)����M��!?  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��L  j�E�P�M�Q�������M��>  ������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��?L  j�U�R�E�P���>����M��6>  ������   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}���K  W�M�Q�U�R���������M�����=  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��K  W�M�Q�U�R����������M�����<  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��TJ  W�M�Q�U�R���4������M����G<  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ���̡���PL���  ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��ZI  j�E�P�M�Q���Y����M��Q;  ������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���H  j�U�R�E�P��������M���:  ������   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��H  j�U�R�E�P���~����M��v:  ������   �
�E�P�у�^��]� ��������U�조��H���   ]��������������U�조��H���   ]�������������̡���H���   �⡰��H���   ��U�조��H���   V�u�R�Ѓ��    ^]�����������U�조��H���   ]��������������U�조��HL�QV�ҋ���u^]á���H�U�Ej R�UP��h  RV�Ѓ���u����Q@�BV�Ѓ�3���^]��������U�조��H�U�E��h  j R�U�� P�ERP�у�]����U�조��H���   ]��������������U�조��H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡���PL�BLQ�Ѓ���������������̡���PL�BPQ�Ѓ����������������U�조��PL�EP�EPQ�JT�у�]� U�조��PL�EPQ��  �у�]� �U�조��PL�EPQ���   �у�]� ̡���PL�BXQ�Ѓ����������������U�조��PL�EP�EP�EPQ�J\�у�]� ������������U���4���SV��HL�QW�ҋ�3ۉ}�;��x  �M���+  ����E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�����   �BSSW���Ѕ���   ����QL�BW�Ћ���;���   ��    ������   �B(���ЍM�Qh�   ���u��
  ������   �M�;���   ������   ���   S��;�tm������   �ȋB<V�Ћ�����   ���   �E�P�у�;�t����B@�HV�у���;��\����}��M��$  �M��+  ��_^[��]� �}�����B@�HW�ы�����   ���   �M�Q�҃��M���#  �M���*  _^3�[��]� �����̡���PL�B`Q�Ѓ���������������̡���PL�BdQ�Ѓ����������������U�조��PL�EPQ�Jh�у�]� ���̡���PL��D  Q�Ѓ������������̡���PL�BlQ�Ѓ����������������U�조��PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh`h@h hR�Q�U R�UR�UR�U���A�$�5���vLRP���   Q�Ѓ�4^]�  ������̡���PL���   Q�Ѓ�������������U�조��PL�EP�EP�EPQ��   �у�]� ���������U�조��PL��H  ]�������������̡���PL��L  ��U�조��PL��P  ]��������������U�조��PL��T  ]��������������U�조��PL��p  ]��������������U�조��PL��t  ]��������������U�조��PL�EP�EP�EP�EP�EPQ���   �у�]� �U�조��PL�EP�EP�EPQ���   �у�]� ���������U�조��PL�EP�EP�EP�EPQ��   �у�]� �����U�조��HL���   ]��������������U�조��HL���   ]��������������U�조��HL���   ]�������������̡���HL��  �⡰��HL��@  ��U�조��PL���  ]��������������U�조��PL���  ]��������������U�조��PL���  ]��������������U��� ���V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\����QLjP���   ���ЋM��U�Rh=���M�}��  ��������   ���   �U�R�Ѓ��M��u��  ��_^��]Ë�����   ���   �E�P�у��M��u���  _�   ^��]����U��� ���V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\����QLjP���   ���ЋM��U�Rh<���M�}���  ��������   ���   �U�R�Ѓ��M��u��L  ��_^��]Ë�����   ���   �E�P�у��M��u��  _�   ^��]����U�조��H��0  ]��������������U��V�u��3�^]ËE�MW�}PQVW��K ����x�V�;�|1�D7� _�F�^]á���H��0  h�QhH  �҃��D7� �F�_^]����������̋A�������������U�조��P8�EPQ�JD�у�]� ���̡���H8�Q<�����U�조��H8�A@V�u�R�Ѓ��    ^]�������������̡���H8�������U�조��H8�AV�u�R�Ѓ��    ^]��������������U�조��P8�EP�EP�EPQ�J�у�]� ������������U�조��P8�EP�EPQ�J�у�]� ����P8�BQ�Ѓ����������������U�조��P8�EPQ�J �у�]� ����U�조��P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U�조��P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�조��P8�EP�EPQ�J(�у�]� U�조��P8�EP�EP�EPQ�J,�у�]� ������������U�조��P8�EP�EP�EPQ�J�у�]� ������������U�조��P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�조��P8�EP�EPQ�J0�у�]� U�조��P8�EP�EP�EPQ�J4�у�]� ������������U�조��P8�EPQ�J8�у�]� ����U�조��H��x  ]��������������U�조��H��|  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H�A,]�����������������U�조��H���  ]��������������U�조��H�QV�uV�ҡ���H�Q8V�҃���^]�����̡���H�Q<�����U�조��H�I@]����������������̡���H�QD����̡���H�QH�����U�조��H�AL]�����������������U�조��H�IP]�����������������U�조��H��<  ]��������������U�조��H��,  ]��������������U�조��H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡���H���   �⡰��H���  ��U�조��H�U�ER�UP�ER�UP���   Rh�2  �Ѓ�]����������������U�조��H�A]�����������������U�조��H��\  ]��������������U�조��H�AT]�����������������U�조��H�AX]�����������������U�조��H�A\]����������������̡���H�Q`�����U�조��H���  ]�������������̡���H�Qd����̡���H�Qh�����U�조��H�Al]�����������������U�조��H�Ap]�����������������U�조��H�At]�����������������U�조��H��D  ]��������������U�조��H��  ]��������������U�조��H�Ix]�����������������U�조��H��@  ]��������������U��V�u���<  ����H�U�A|VR�Ѓ���^]���������U�조��H���   ]��������������U�조��H��h  ]��������������U�조��H��d  ]��������������U�조��H���  ]�������������̡���H���   ��U�조��H��l  ]��������������U�조��H��   ]��������������U�조��H��  ]��������������U��V�u����  ����H���   V�҃���^]���������̡���H��`  ��U�조��H��  ]��������������U�조��H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U�조��H���  ]��������������U��U�E����H�E���   R���\$�E�$P�у�]�U�조��H���   ]��������������U�조��H���   ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���   ]��������������U�조��H���   ]��������������U�조��H���   ]��������������U�조��H���   ]��������������U�조��H���   ]��������������U�조��H���   ]��������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�조��H��8  ]��������������U��V�u(V�u$�E�@����R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@����R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�조��P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�조��P0�EP�EP�EP�EPQ���   �у�]� ����̡���P0���   Q�Ѓ�������������U�조��P0�EP�EPQ���   �у�]� �������������U�조��P0�EP�EP�EP�EPQ���   �у�]� ����̡���P0���   Q�Ѓ������������̡���H0���   ��U�조��H0���   V�u�R�Ѓ��    ^]�����������U�조��H��H  ]��������������U�조��H��T  ]�������������̡���H��p  �⡰��H���  ��U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ������   �Qj PV�ҡ�����   ��U�R�Ѓ� ��^��]��������U���4VhLGOg�M��l  ����Q��X  3�VP�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�у� �M��R  ������   �PT�M�Q�҃���u'�u����  ������   ��U�R�Ѓ���^��]Ë�����   �JT�E�P�ыu��P����  ������   ��M�Q�҃���^��]���������������U�조��H��  ]��������������U�조��H��\  ]��������������U�조��H�U��t  ��V�uVR�E�P�у����4  �M���3  ��^��]�����U�조��H�U���  ��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]����������������U�조��H�U���  ��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]����������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H�U�E��VWj R�UP�ERP��t  �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�(_��^��]��U�조��H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у�$��^��]���U�조��H��8  ]��������������U���  ��3ŉE��M�EPQ������h   R�8 ����x	=�  |#�����H��0  h�QhH  �҃��E� ����H��4  ������Rh�Q�ЋM�3̓��C�  ��]�������U��E�M�UPQRhR�W�������H��0  h�Qh�  �҃�]���������U�조��H��  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]����U�조��H��  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]����U�조��H��p  ��4�҅���   h���M���  ����P�E�R4Ph���M��ҡ���P�E�R4Ph���M��ҡ���H��X  j �U�R�E�hicMCP�ы���E�    �E�    ���   j P�A�U�R�Ћ�����   �
�E�P�ы�����   ��M�Q�҃�$�M��[  ��]��������U�조��H��p  ��4V�҅�u����H�u�QV�҃���^��]�Wh!���M���  ����P�E�R4Ph!���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �PH�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ�����   ��U�R�Ѓ�4�M��M  _��^��]������U�조��H��p  ��4V�҅�u����H�u�QV�҃���^��]�Wh����M��  ����P�E�R4Ph����M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �PH�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ�����   ��U�R�Ѓ�4�M��=  _��^��]������U�조��H��p  ��4�҅�u��]�Vh#���M���  ����P�E�R4Ph#���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �P8�M�Q�ҋ�����   ��U�R�Ѓ�(�M��e  ��^��]���������������U�조��H��p  ��4�҅�u��]�Vhs���M���  ����P�E�R4Phs���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �P8�M�Q�ҋ�����   ��U�R�Ѓ�(�M��  ��^��]���������������U�조��H���  ]��������������U�조��H��@  ]��������������U�조��H���  ]��������������U��V�u���t����QP��D  �Ѓ��    ^]������U�조��H��H  ]��������������U�조��H��L  ]��������������U�조��H��P  ]��������������U�조��H��T  ]��������������U�조��H��X  ]��������������U�조��H��\  ]�������������̡���H��d  ��U�조��H��h  ]��������������U�조��H��l  ]�������������̡���H���  ��U�조��H�U���  ��VR�E�P�ыu��P���s	  �M��	  ��^��]�����U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H��l  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H��$  ]��������������U�조��H��(  ]��������������U�조��H��,  ]�������������̡���H��0  �⡰��H��<  ��U�조��H���  ]�������������̡���H���  ��U�조��H���  ]��������������U��Q�Mj �  �E���tP�����E�P��M������]������U�조��H��  ]�������������̡���H��P  ��U�조��H��`  ]�������������̡�����   ���   ��Q��Y��������U�조��H�A�U��� R�Ћ���Q�Jj j��E�h$RP�ы���B�P�M�Q�ҡ���H�I�U�R�E�P�ы���B�P<�� �M��ҋ���Q�M�RLj�j�QP�M��ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�҃���]��������������U�조��P�B<V���Ћ���Q�M�RLj�j�QP���ҋ�^]� �������������U�조��H�QV�uV�ҡ���H�U�AVR�Ћ���Q�B<�����Ћ���Q�M�RLj�j�QP���ҋ�^]��������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���I  �����   �ESP�M��X#  ����Q�J�E�P�ы���B�Pj j��M�h$QQ�҃��E�P�M��#  j j��M�Q�U�R��d���P�8  ��P�M�Q�'  ��P�U�R�
'  ���P�J  ���M����Q#  �M��I#  ��d����>#  �M��6#  ����H�A�U�R�Ѓ��M��#  ��[t	V�H  ����^��]� ���U��EVP���aS  �����^]� �����Q�H  Y���������U��E�M�U�H4�M�P �U��M�@p} �@80.�@<p.�@@�.�@D�-�@H�.�@L@.�@P .�@lP.�@X�.�@\.�@`�.�@d`.�@T�.�@h�.�@p�-�@t .�P0�H(�@,    ]��������������U���   h�   ��`���j P���  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj������8��]��������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,����������̡�����   �BQ�Ѓ������������̡�����   �BXQ�Ѓ�������������U�조����   �EPQ�J`�у�]� �U�조��P���   ]�������������̡���P�B�����U�조��P�Rt]�����������������U�조��P�Rl]����������������̡���P�BVj j����Ћ�^���������U�조��P�E�RVj P���ҋ�^]� U�조��P�E�RVPj����ҋ�^]� ����P�B�����U�조��P���   Vj ��Mj V�Ћ�^]� �����������U�조��P�EPQ�J�у�]� ����U�조��P�EPQ�J�у����@]� ���������������U�조��P�E�RtP�ҋ�����   P�BX�Ѓ�]� ���U�조��P�E�Rlh#  P�EP��]� ���������������U�조��P�E�RlhF  P�EP��]� ���������������U�조��P�E�RtP�ҋ�����   �M�R`QP�҃�]� ���������������U�조��P���   ]��������������U�조��P�E���   P�҅�u]� ������   P�B�Ѓ�]� �������̋��     �@    á���PD�BQ�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�BQ�Ѓ����������������U�조��PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U�조��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�조��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�조��PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U�조��PX�EPQ�J�у�]� ����U�조��PX�EPQ�J�у�]� ����U�조��PX�EPQ�J�у�]� ����U�조��PX�EPQ�J�у�]� ����U�조��PX�EPQ�J$�у�]� ����U�조��PX�EPQ�J �у�]� ����U�조��PD�EP�EPQ�J�у�]� U�조��HD�U�j R�Ѓ�]�������U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��HD�	]��U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��HD�U�j R�Ѓ�]�������U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��U�HD�Rh2  �Ѓ�]����U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��U�HD�RhO  �Ѓ�]����U�조��H@�AV�u�R�Ѓ��    ^]��������������U�조��U�HD�Rh'  �Ѓ�]����U�조��H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h�  �҃�����������U�조��H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h:  �҃�����������U�조��H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E�������   �R�E�Pj�����#E���]�̡���HD�j h�F �҃�����������U�조��H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h�_ �҃�����������U�조��H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E�����E�    ���   �R�E�Pj������؋�]� ̡���PD�B$Q�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ����������������h��PhD � O  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h��jhD �LN  ����t
�@��t]��3�]��������Vh��j\hD ���N  ����t�@\��tV�Ѓ���^�����Vh��j`hD ����M  ����t�@`��tV�Ѓ�^�������U��Vh��jdhD ���M  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh��jhhD ���yM  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh��jlhD ���<M  ����t�@l��tV�Ѓ�^�������U��Vh��h�   hD ���M  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh��h�   hD ���L  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh��jphD ���iL  ����t�@p��t�MQV�Ѓ�^]� ���^]� ��U��Vh��jxhD ���)L  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh��j|hD ����K  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh��j|hD ���K  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vh��h�   hD ���SK  ����t=���   ��t3�MQ�U�VR��h��j`hD �&K  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������h��jhD ��J  ����t	�@��t��3��������������U��V�u�> t+h��jhD �J  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h��jhD �aJ  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh��jhD ���J  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh��jhD ����I  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh��j hD ���I  ����t�@ ��tV�Ѓ�^�3�^���Vh��j$hD ���lI  ����t�@$��tV�Ѓ�^�3�^���U��Vh��j(hD ���9I  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh��j,hD ����H  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh��j(hD ���H  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh��j4hD ���\H  ����t�@4��tV�Ѓ�^�3�^���U��Vh��j8hD ���)H  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh��j<hD ����G  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh��jDhD ���G  ����t�@D��tV�Ѓ�^�3�^���U��Vh��jHhD ���iG  ����t�M�PHQV�҃�^]� U��Vh��jLhD ���9G  ����u^]� �M�PLQV�҃�^]� �����������U��Vh��jPhD ����F  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh��jThD ���F  ����u^Ë@TV�Ѓ�^���������U��Vh��jXhD ���F  ����t�M�PXQV�҃�^]� U��Vh��h�   hD ���VF  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh��h�   hD ���F  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh��h�   hD ���E  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���vE  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���6E  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ����D  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh��h�   hD �D  ����u����H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]��U��Vh��h�   hD ���&D  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   hD ����C  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   hD ���C  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   hD ���VC  ����t���   ��t�MQ����^]� 3�^]� �Vh��h�   hD ���C  ����t���   ��t��^��3�^����������������U��Vh��h�   hD ����B  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   hD ���B  ����t���   ��t�MQ����^]� ��������U��Vh��h�   hD ���FB  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh��h�   hD ����A  ����t���   ��t��^��3�^����������������VW��3����$    �h��jphD �A  ����t�@p��t	VW�Ѓ������8 tF��_��^�������U��SW��3�V��    h��jphD �_A  ����t�@p��t	WS�Ѓ������8 tqh��jphD �-A  ����t�@p��t�MWQ�Ѓ�������h��jphD ��@  ����t�@p��t	WS�Ѓ�����V���������tG�]����E^��t�8��~=h��jphD �@  ����t�@p��t	WS�Ѓ������8 u_�   []� _3�[]� ����������U��Vh��j\hD ���Y@  ����t3�@\��t,V��h��jxhD �7@  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh��j\hD ����?  ����t3�@\��t,V��h��jdhD ��?  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh��j\hD ���?  ����tG�@\��t@V�ЋEh��jdhD �E��E�    �E�    �`?  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��j\hD ���?  ����t\�@\��tUV��h��jdhD ��>  ����t�@d��t
�MQV�Ѓ�h��jhhD ��>  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh��j\hD ���>  ������   �@\��t~V��h��jdhD �c>  ����t�@d��t
�MQV�Ѓ�h��jhhD �:>  ����t�@h��t
�URV�Ѓ�h��jhhD �>  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh��jthD ����=  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h��j`hD �=  ����th�@`��ta�M�Q�Ѓ���^��]� h��j\hD �m=  �u����t4�@\��t-V��h��jdhD �H=  ����t�@d��th��V�Ѓ���^��]� ������U���Vh��h�   hD �=  ����tU���   ��tK�M�UQR�M�Q�Ћu��P���h���h��j`hD ��<  ����te�@`��t^�U�R�Ѓ���^��]�h��j\hD �<  �u����t3�@\��t,V��h��jxhD �s<  ����t�@x��t
�MVQ�Ѓ���^��]�����U���Vh��h�   hD ���3<  ����tR���   ��tH�MQ�U�R���ЋuP������h��j`hD ��;  ����t|�@`��tu�M�Q�Ѓ���^��]� h��j\hD �E�    �E�    �E�    �;  �u����t3�@\��t,V��h��jdhD �;  ����t�@d��t
�U�RV�Ѓ���^��]� ��������������U�조��UV��H�AVR�Ѓ���^]� ��������������U�조��P�Rd]�����������������U�조��P�Rh]�����������������U�조��P�EP�EP�EPQ�J�у�]� �����������̡��V��H�QV�ҡ���H$�QDV�҃���^�����������U�조�V��H�QV�ҡ���H$�QDV�ҡ���U�H$�AdRV�Ѓ���^]� ��U�조�V��H�QV�ҡ���H$�QDV�ҡ���U�H$�ARV�Ѓ���^]� ��U�조�V��H�QV�ҡ���H$�QDV�ҡ���H$�U�ALVR�Ѓ���^]� �̡��V��H$�QHV�ҡ���H�QV�҃�^�������������U�조��P$�EPQ�JL�у�]� ����U�조��P$�R]�����������������U�조��P$�Rl]����������������̡���P$�Bp����̡���P$�BQ�Ѓ����������������U�조��P$��VWQ�J�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]� ���U�조��P$�EPQ�J�у�]� ����U�조��P$��VWQ�J �E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]� ���U�조��P$��VWQ�J$�E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]� ���U���,VW�E�P�o�������Q$�JP�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у� _��^��]� �����̡���P$�B(Q��Yá���P$�BhQ��Y�U�조��P$�EPQ�J,�у�]� ����U�조��P$�EPQ�J0�у�]� ����U�조��P$�EPQ�J4�у�]� ����U�조��P$�EPQ�J8�у�]� ����U�조��UV��H$�ALVR�Ѓ���^]� ��������������U�조��H�QV�uV�ҡ���H$�QDV�ҡ���H$�U�ALVR�Ћ���E�Q$�J@PV�у���^]�U�조��UV��H$�A@RV�Ѓ���^]� ��������������U�조��P$�EPQ�J<�у�]� ����U�조��P$�EPQ�J<�у����@]� ���������������U�조��P$�EP�EPQ�JP�у�]� U�조��P$�EPQ�JT�у�]� ���̡���H$�QX�����U�조��H$�A\]�����������������U�조��P$�EP�EP�EPQ�J`�у�]� �����������̡���H(�������U�조��H(�AV�u�R�Ѓ��    ^]��������������U�조��P(�R]����������������̡���P(�B�����U�조��P(�R]�����������������U�조��P(�R]�����������������U�조��P(�R ]�����������������U�조��P(�E�RjP�EP��]� ��U�조��P(�E�R$P�EP�EP��]� ����P(�B(����̡���P(�B,����̡���P(�B0�����U�조��P(�R4]�����������������U�조��P(�RX]�����������������U�조��P(�R\]�����������������U�조��P(�R`]�����������������U�조��P(�Rd]�����������������U�조��P(�Rh]�����������������U�조��P(�Rl]�����������������U�조��P(�Rx]�����������������U�조��P(���   ]��������������U�조��P(�Rt]�����������������U�조��P(�Rp]�����������������U�조��P(�BpVW�}W���Ѕ�t:����Q(�Rp�GP���҅�t"����P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U�조��P(�BtVW�}W���Ѕ�t:����Q(�Rt�GP���҅�t"����P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U�조��P(�BpSVW�}W���Ѕ���   ����Q(�Rp�GP���҅���   ����P(�Rp�GP���҅�tp����P(�Bp�_S���Ѕ�tY����Q(�Rp�CP���҅�tA����P(�Bp��S���Ѕ�t*�OQ��������t��$W��������t_^�   []� _^3�[]� ���U�조��P(�BtSVW�}W���Ѕ���   ����Q(�Rt�GP���҅���   ����P(�Rt�GP���҅�tp����P(�Bt�_S���Ѕ�tY����Q(�Rt�CP���҅�tA����P(�Bt��S���Ѕ�t*�O0Q���+�����t��HW��������t_^�   []� _^3�[]� ���U�������E�    �E�    �P(�RhV�E�P���҅���   �E���uG����H�A�U�R�Ћ���Q�E�RP�M�Q�ҡ���H�A�U�R�Ѓ��   ^��]� ����Qh(Rhe  P���   �Ћ�����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�����3�^��]� ����E��Q�M�j HP�EQ�JP�эU�R�������   ^��]� �����U�조���V��H�A�U�R�Ѓ��M�Q������^��u����B�P�M�Q�҃�3���]� ����H$�E�I�U�RP�ы���B�P�M�Q�҃��   ��]� �U��Q����P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U�조��P(�R8]�����������������U�조��P(�R<]�����������������U�조��P(�R@]�����������������U�조��P(�RD]�����������������U�조��P(�RH]�����������������U�조��P(�E�R|P�EP��]� ����U�조��P(�RL]�����������������U�조��E�P(�BT���$��]� ���U�조��E�P(�BPQ�$��]� ����̡���H(�Q�����U�조��H(�AV�u�R�Ѓ��    ^]��������������U�조��P(���   ]��������������U�조��H(�A]����������������̡���H,�Q,����̡���P,�B4�����U�조��H,�A0V�u�R�Ѓ��    ^]�������������̡���P,�B8�����U�조��P,�R<��VW�E�P�ҋu������H�QV�ҡ���H$�QDV�ҡ���H$�QLVW�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у�_��^��]� �������U�조��P,�E�R@��VWP�E�P�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ��̡���H,�j j �҃��������������U�조��P,�EP�EPQ�J�у�]� U�조��H,�AV�u�R�Ѓ��    ^]�������������̡���P,�B����̡���P,�B����̡���P,�B����̡���P,�B ����̡���P,�B$����̡���P,�B(�����U�조��P,�R]�����������������U�조��P,�R��VW�E�P�ҋu������H�QV�ҡ���H$�QDV�ҡ���H$�QLVW�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у�_��^��]� �������U�조��H��D  ]��������������U�조��H��H  ]��������������U�조��H��L  ]��������������U�조��H�I]�����������������U�조��H�A]�����������������U�조��H�I]�����������������U�조��H�A]�����������������U�조��H�I]�����������������U�조��H���  ]��������������U�조��H�A]�����������������U���V�u�E�P����������Q$�J�E�P�у���u-����B$�PH�M�Q�ҡ���H�A�U�R�Ѓ�3�^��]Ë���Q�J�E�jP�у���u=�U�R��������u-����H$�AH�U�R�Ћ���Q�J�E�P�у�3�^��]Ë���B�HjV�у���u����B�HV�у����I�������Q$�JH�E�P�ы���B�P�M�Q�҃��   ^��]�����������U�조��H�A ]�����������������U�조��H�I(]�����������������U�조��H��  ]��������������U�조��H��   ]��������������U�조��H��  ]��������������U�조��H��  ]��������������U�조��H�A$��V�U�WR�Ћ���Q�u���BV�Ћ���Q$�BDV�Ћ���Q$�BLVW�Ћ���Q$�JH�E�P�ы���B�P�M�Q�҃�_��^��]������U�조��H���  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q$�BDV�Ћ���Q$�BLVW�Ћ���Q$�JH�E�P�ы���B�P�M�Q�҃�_��^��]���U�조��H���  ]��������������U���<���SVW�E�    ��t�E�P�   �������/����Q�J�E�P�   �ы���B$�PD�M�Q�҃��}ࡰ��H�u�QV�ҡ���H$�QDV�ҡ���H$�QLVW�҃���t)����H$�AH�U�R����Ћ���Q�J�E�P�у���t&����B$�PH�M�Q�ҡ���H�A�U�R�Ѓ�_��^[��]���U�조��H�U���  ��VWR�E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]��������������U�조��H���  ]�������������̡���H���   ��U�조��H���   V�uV�҃��    ^]�������������U�조��P�]�⡰��P�B����̡���P���   ��U�조��P�R`]�����������������U�조��P�Rd]�����������������U�조��P�Rh]�����������������U�조��P�Rl]�����������������U�조��P�Rp]�����������������U�조��P�Rt]�����������������U�조��P���   ]��������������U�조��P��  ]��������������U�조��P�Rx]�����������������U�조��P���   ]��������������U�조��P�R|]�����������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P�EPQ��  �у�]� �U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U��E��t ����R P�B$Q�Ѓ���t	�   ]� 3�]� U�조��P �E�RLQ�MPQ�҃�]� U��E��u]� ����R P�B(Q�Ѓ��   ]� ������U�조��P�R]�����������������U�조��P�R]�����������������U�조��P�R]�����������������U�조��P�R]�����������������U�조��P�R]�����������������U�조��P�R]�����������������U�조��P�E�R\P�EP��]� ����U�조��P�E��  P�EP��]� �U�조��E�P�B ���$��]� ���U�조��E�P�B$Q�$��]� �����U�조��E�P�B(���$��]� ���U�조��P�R,]�����������������U�조��P�R0]�����������������U�조��P�R4]�����������������U�조��P�R8]�����������������U�조��P�R<]�����������������U�조��P�R@]�����������������U�조��P�RD]�����������������U�조��P�RH]�����������������U�조��P�RL]�����������������U�조��P�RP]�����������������U�조��P���   ]��������������U�조��P�RT]�����������������U�조��P�EPQ��  �у�]� �U�조��P���   ]��������������U�조��P���   ]��������������U�조��P�RX]����������������̡���P���   ��U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]��������������U�조��P���   ]�������������̡���P���   ��U�조��P���   ]�������������̡���P���   �ࡰ��P���   �ࡰ��P���   ��U�조��H���   ]��������������U�조��H��   ]��������������U�조��H�U�E��VWRP���  �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]������������U�조��H���  ]��������������U�조��P(�BPVW�}�Q�]���E�$�Ѕ�tM����G�Q(�]�E�BPQ���$�Ѕ�t,����G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U�조��P(�BTVW�}����$���Ѕ�tE����G�Q(�BT�����$�Ѕ�t(����G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U�조��P(�BTVW�}����$���Ѕ�tr����G�Q(�BT�����$�Ѕ�tU����G�Q(�BT�����$�Ѕ�t8�OQ���������t)�W0R��������t��HW��������t_�   ^]� _3�^]� ���U�조��P(�} �R8����P��]� �U�조��P�BdS�]VW��j ���Ћ���Qh(R�p���   h�  V�Ћ�����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ���Q(�BHV���Ѕ�t ����Q(�E�R VP���҅�t�   �3��EP�r����_��^[]� ������U�조��U�� V��H$�IWR�E�P�ы�����B�P�M�Q�ҡ���H�A�U�RW�Ћ���Q�J�E�P�у��U�R�����������H�A�U�R�Ѓ�_��^��]� �����������U�조��P|�EP�EPQ�J8�у�]� U�조����   �BXQ�Ѓ���u]� ����Q|�M�RQ�MQP�҃�]� ���U�조����   �BXQ�Ѓ���u]� ����Q|�M�R8Q�MQP�҃�]� ���U��EV��j �����Qj j P�B�ЉF����^]� ��̡��Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ����Q�MP�EP�Q�JP�у��F�   ^]� ����U��E#E]�����̋�3ɉ�H�H�H�H�H�����������V���h���3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX��^��̡���P�BQ�Ѓ���������������̡���P�BQ�Ѓ���������������̡���H���   ��U�조��H���   V�u�R�Ѓ��    ^]����������̡���P���   Q�Ѓ�������������U�조��P�EPQ���   �у�]� ̡���H�������U�조��H�AV�u�R�Ѓ��    ^]��������������U�조��H�AV�u�R�Ѓ��    ^]��������������U�조��P��Vh�  Q���   �E�P�ы�����   �Q8P�ҋ�����   ��U�R�Ѓ���^��]��������������̡���P�BQ�Ѓ����������������U�조��P�EPQ�J\�у�]� ����U�조��P�EP�EP�EP�EP�EPQ���   �у�]� �U�조��P�EP�EP�EP�EPQ�JX�у�]� �������̡���P�B Q��Y�U�조��P�EP�EP�EP�EPQ���   �у�]� �����U�조��P�EP�EP�EPQ�J�у�]� ������������U�조��H��   ]��������������U�조��P�R$]�����������������U�조��P��x  ]�������������̡���P��|  ��U�조��P�EP�EP�EP�EPQ�J(�у�]� ��������U�조��P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U�조��P�EP�EP�EP�EPQ�J,�у�]� ��������U�조�V��H�QWV�ҍx�����H�QV�ҋ���Q�M�R4Q�MQ�MQWHPj j V�҃�(_^]� ���������������U�조��P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U�조��P�EP�EPQ�J@�у�]� U�조��P�EPQ�JD�у�]� ���̡���P�BLQ�Ѓ���������������̡���P�BLQ�Ѓ���������������̡���P�BPQ�Ѓ����������������U�조��P�EPQ�JT�у�]� ����U�조��P�EPQ�JT�у�]� ����U�조��P�EP�EPQ���   �у�]� �������������U�조��P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у� ��^��]� ������̡���P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡���H�������U�조��H�AV�u�R�Ѓ��    ^]��������������U�조��P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�조��P�EPQ�J�у�]� ���̡���P�BQ��Y�U�조��P�EP�EPQ�J�у�]� U��VW�������M�U�x@�EPQR�������H ���_^]� �U��VW������M�U�xD�EPQR������H ���_^]� �V������xH u3�^�W���v���΍xH�l���H �_^�����U��V���U���xL u3�^]� W���@���M�U�xL�EPQR���*���H ���_^]� �������������U��V������xP u���^]� W���� ���M�U�xP�EP�EQRP���� ���H ���_^]� ��������U��V��� ���xT u���^]� W��� ���M�xT�EPQ��� ���H ���_^]� U��V���u ���xX u���^]� W���_ ���xX�EP���Q ���H ���_^]� ����U���S�]VW���t.�M��V������ ���xL�E�P��� ���H ��ҍM�萲���}��tZ����H�A�U�R�Ћ���Q�J�E�WP�ы���B�P�M�Q�҃��������@@��t����QWP�B�Ѓ�_^[��]� ������U��V�������x` u
� }  ^]� W���m����x`�EP���_����H ���_^]� ��U��VW���D����xH�EP���6����H ���_^]� ���������U��SVW�������x` u� }  �#��������x`�E���P��������H ��ҋ�����H�]�QS�҃�;�A����H�QS�҃�;�,�������M�U�xD�EPQSR�������H ���_^[]� _^�����[]� ��������������U��V���e����xP u
�����^]� W���M����M�U�xP�EP�EQ�MR�UPQR���+����H ���_^]� ��������������U��V�������xT u
�����^]� W��������M�xT�EPQ��������H ���_^]� ��������������U��V�������xX tW�������xX�EP�������H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u���>  ����t.�E�;�t'����J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡���H��   ��U�조��H��$  V�u�R�Ѓ��    ^]�����������U�조��UV��H��(  VR�Ѓ���^]� �����������U�조��P�EQ��,  P�у�]� �U�조��P�EQ��,  P�у����@]� �����������̡���H��0  �⡰��H��4  �⡰��H��p  �⡰��H��t  ��U��E��t�@�3�����RP��8  Q�Ѓ�]� �����U�조��P�EPQ��<  �у�]� �U�조��P�EP�EP�EPQ��@  �у�]� ���������U�조��P�EP�EPQ��D  �у�]� �������������U�조��P�EPQ��H  �у�]� �U�조��P�E��L  ��VWPQ�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ��������������̡���P��T  Q�Ѓ�������������U�조��P�EPQ��l  �у�]� ̡���P��P  Q�Ѓ�������������U�조��P�EPQ��X  �у�]� ̡���H��\  ��U�조��H��`  V�u�R�Ѓ��    ^]�����������U�조��P�EP�EP�EP�EP�EPQ��d  �у�]� �U�조��P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���O�������3��G �G$�G(�G,�G0�G4�G8�G<�G@�GD�GH�GL�GP�GT�GX�G\�_p��G`�Gd�Gh�Gx�����G|   ��_^����������������V��W�>��t7���/����xP t$S���!���j j �XPj�FP�������H ���[�    �~` t����H�V`�AR�Ѓ��F`    _^������������U��SV��Fx����Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�$�������u#���h\R����H��0  h  �҃��E�~P�������j j jW�����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ����Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��QV��~d tg�E;Fxt_�N`W�>�M����{����xP u����(S���h����UR�XP�E�Pj�NQ���P����H ���[�F|_��u�E�Fx�E��t�    �F`^��]� �M�Fx������t�3�^��]� ���������U��QVW�}����;  ����H�QhV�҃������u"�H��0  h\Rh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���?9  �EF;u�|�UR�m�����_�   ^��]� �������������U��QVW�}�����:  ����H�QhV�҃������u"�H��0  h\Rh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'������QP�Bh�Ѓ���t�M��R���\8  F;u�|ʍEP������_�   ^��]� �������������h\Rh�   h��h�   �W�������t������3��������V��������N^�/������������������U��VW�}�7��t�������N����V�=������    _^]�����������������U��]�7  ��������{9  �����������U��]�w7  ��������[9  �����������U��V���E����N�����Et	V���������^]� �������U��E�M�UP��P�EjP������]��������������̸   �����������U��V�u��t���u6�EjP��������u3�^]Ë�������t���t��U3�;P��I#�^]������̡���H\�������U�조��H\�AV�u�R�Ѓ��    ^]�������������̡���P\�BQ�Ѓ���������������̡���P\�BQ�Ѓ����������������U�조��P\�EPQ�J�у�]� ����U�조��P\�EP�EPQ�J�у�]� U�조��P\�EPQ�J�у�]� ���̡���P\�BQ�Ѓ����������������U�조��P\�EPQ�J �у�]� ����U�조��P\�EP�EPQ�J$�у�]� U�조��P\�EP�EP�EP�EPQ�J`�у�]� ��������U�조��P\�EPQ�J0�у�]� ����U�조��P\�EPQ�J@�у�]� ����U�조��P\�EPQ�JD�у�]� ����U�조��P\�EPQ�JH�у�]� ���̡���P\�B4Q�Ѓ����������������U�조��P\�EP�EPQ�J8�у�]� U�조��P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu���������H\�QV�҃���S������3���~B��I ����H\�U�R�U��EP�A`h���VR�ЋM��Q���S����U�R���H���F;�|�_^[��]� ����������U���VW�}�E��P���x����}� ��   ����Q\�BV�Ѓ��M�Q���Q����E���t]S3ۅ�~H�I �UR���5����E�P���*����E;E�!������Q\P�BV�ЋE@���E;E�~�C;]�|�[_�   ^��]� _�   ^��]� U��M�EV�uIH��tS�Y�PA@N��u�[^]� �������U��M�EV�u������t!W���    �Pf�y����Nf�8f�u�_^]� ���U��M�EV�u������tW���    �y�P����N�8�u�_^]� �������U��� �E�M���  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��4�E��}���t�u+��\�P@�M���u�EH�E����   )}��u��	;]��u��s���u�]�;]}�M��>P�E�V�Ѕ�y�u�C�]�M��E��VP�҅��d����F��}��t�M�+���I ��P@�M��T�u�]��;]~��/���_^[��]� ������U���(W�}�����E�E�M���/  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��
�U���$    ��~�M�M�J)}��U��G�M�E��M��t'�M�+����$    ��pf�\���M�f�f�4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��H����}�F���t!�M�+ȍI �Pf���Of�f�T�u�]��}�;E�~����	���^[_��]� ����������U���(W�}�����E�E�M���  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��9�M�E��M��t�M�+ȋ\�p���M��4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��W����}�F���t�M�+Ȑ��P��O��T�u�]��}�;E~��"���^[_��]� ��U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   xO�E�   �}��}_^3�[��]� �}}���E������uu��VP�҅�tyO�}�G�}��E9E�~�_^3�[��]� ��~3�E���]��]�E����E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   y�M_^�    3�[��]� �O�3��E�   �M��} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�ty�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U���E]鴎  ����U���E��]�������U���E����P�X]� �����������̋�� �����������U����M�� ��A�@�X�A�@�X]� ������������U��U�M�B�I�E�A�J����A�
�B�	���X�B�	��I���X]�����U��V�u�F��F�����������������܍  ��������������D�Ez��^��P�X]��������������N�X�N^�X]���������������U��M�U��"�E��A�b�X�A�b�X]����������������P�P�P�P �P(�P0�P8�P@�PH�PP�PX����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX�������̋�� �����������U��M�U�A�
�E��A0�J���AH�J����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X]����U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH������������Dz�u�؋��������^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]����̋%    ��������̋�   @t���Ã����������������������P�P�P�P �X(��R�@0    ��������X�X��R�������X�X �X(�����������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A�A �A�A(��P����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E������X�X]� ̋�3ɉ�H�H�H�V��V�g����FP�^���3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}��+	  S�]����  ��؋���M�U��>���U�@�U���� �U��@�@�B�@�������@���@�   ���]��E��U�;���  �w�����  �w�������F�ݍB��   �U����������������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]����]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]��]��U���E��U��R�э����N�B���B�P���R���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]�����B���B���U����E��������]��E����E����������E������E��E��U����E��]����E��U��E��U��P����E�̋U���������������;���   �ލ���+�������̋�@�������O�]��@���]��@���U������M������]��E��E����E������E����������E��E��U����E��]����E��U��E��E��U�u�����������������������[�[�E��������������L�  ��������������Dz���������E��-������������������M����M��E��������������������[H���[P�[X�E����E���������zu������������zh�����CP���CX���CH���CX�������cH���[���[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@��   ������������z]�CX���CP�����cH�CH���CP�������[�[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@�]�CP���CX�����CH���CX�����cP���[0���[8�[@�C8�KX�C@�KP���CH�K@�C0�KX���C0�KP�C8�KH�����[�[ �[(��$���SQ�����E��U�   �����}��M������3�3��u��u���|)�A�����B�4�u�0u��u�p��J�u�u�U�E;�}�Q���E���u��U��1���@���K�I�E    ��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]�� �K��C0�H���@�KH��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���U����n  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������]��E�E����]���E����]��E��M����@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������U��E��]��E��U������������������9M|��[��_��^���؋�]� ���������ʋE�����׋��@�E�Ѝ��K��C0�H���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���CX�H�E@�E���]����E��������������������M����������]��E��E�;��T�����[������_��^��]� �h��Ph_� �������������������h��jh_� �_�������uË@����U��V�u�> t/h��jh_� �3�������t��U�M�@R�Ѓ��    ^]���U��Vh��jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh��jh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh��jh_� ���y�������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jh_� ���)�������t�@��t�MQ����^]� 3�^]� �������U��Vh��j h_� �����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh��j$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh��j(h_� ���l�������t�@(��t��^��3�^������Vh��j,h_� ���<�������t�@,��t��^��3�^������U��Vh��j0h_� ���	�������t�@0��t�MQ����^]� 3�^]� �������U��Vh��j4h_� �����������t�@4��t�M�UQR����^]� ���^]� ��Vh��j8h_� ����������t�@8��t��^��3�^������U��Vh��j<h_� ���Y�������t�@<��t�MQ����^]� ��������������U��Vh��j@h_� ����������t�@@��t�MQ����^]� ��������������U��Vh��jDh_� �����������t�@D��t�MQ����^]� 3�^]� �������U��Vh��jHh_� ����������t�@H��t�MQ����^]� ��������������Vh��jLh_� ���\�������t�@L��t��^��3�^������Vh��jPh_� ���,�������t�@P��t��^��3�^������Vh��jTh_� �����������t�@T��t��^��^��������Vh��jXh_� �����������t�@X��t��^��^��������Vh��j\h_� ����������t�@\��t��^��^��������U��Vh��j`h_� ���i�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh��jdh_� ���)�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh��jhh_� �����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh��jlh_� ����������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jph_� ���I�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh��jth_� ���	�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh��jxh_� �����������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh��j|h_� ����������t�@|��t�MQ����^]� 3�^]� �������U��Vh��h�   h_� ���F�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh��h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh��h�   h_� ���6�������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h_� �����������t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   h_� ����������t���   ��t�MQ����^]� ��������U��Vh��h�   h_� ���f�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h_� ����������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E����������M������U�_��^�U�[���U������������������������'t  ��������������D�Ez����P�X��]� �������E�����E����X�M��X��]� ��U���@��R�A���E�    �����]��]��]���R�������]��]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�1����F�@��R�M������~���Q�M������v;�t�v��P�M�������M����M��M�u�_^[�M�UQR�M�������]� �Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��x+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~!V�1�d$ ���   @u	�����t@��Ju�^�����̋QV3���~�	�d$ ����ШtF��Ju��^�����������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%����E���;�}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�(��E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��±ر��������U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP����3����F�F^��U��SV��WV�����^S�����E3����~�~;�t_����Q���   h�R��jIP�у��;�t9�}��t;����B���   h�R��    jNQ�҃����uV������_^3�[]� �E�~_�F^�   []� ����������U��V��WV������FP������}���F    �F    ����   �? ��   �G����   ����Q���  h�R��jlP�у����t>� t@�G��t9����Jh�R��    ���  jqR�Ѓ��F��u�������_3�^]� �O��N�G�F��    ���t��t��tQPR�Sd  ���F��t�VP��RP�GP�  ��_�   ^]� ��������U��SV��WV������~W�����3����F�F9E�  �];���   ����Qh�R��    h�   P���  �Ѓ����t@�} tN�]��tD����Q���  h�R��    h�   P�у����u�������_^3�[]� �^�]�0�]�F   ����B���  h�Rh�   j�у����t���^��t��    ��t�UQRP�c  ���E��t!�N�?�W�QWP�R  ��_^�   []� ��_^�   []� ���U��Q�A�E� ��~JS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U���Ou�_^[�E��Ћ�]� �����������U��S�]V��3�W�~���F�F�CV;C��   ����W�����3��F�F����Q���   h�RjIj�Ѓ������   ����Q���   h�RjNj�Ѓ����uV覿����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �`���W�Z���3��F�F����B���   h�RjIj�у����t[����B���   h�RjNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�`  ��]�����������̋�   @u
���ȃ��u3�ø   �����U�조��H�U�I(��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]���U�조��E�H�U �E��VWR�UP�ERP�A$���U��$R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�,_��^��]��������������U��Q����P�E�RdWP�M��ҋ���u_��]� ����H���   SVh�R�_j	S�ҋ�����u	^[_��]� ����P�E�M��RhPSV���> ��^[_��]� ������U�����3ŉE�S�]VW�}f�E�0x�   �   ��$    �ǋ���$<
}0�7�D�B��y����D� �Q�BS�Ћ���Q�Jj j��E�PS�ыM���_^��3�[��c  ��]����U���0V�uW�}����  ��   @�  ����H�A�U�R�Ћ���Q�Jj j��E�h0SP�ы���B�P$����j0��j �}�ujj �m���M��(S�$Q�ҋ���H�A�U�R�Ћ���Q�J�E�PV�ы���B�P�M�Q�ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�B<��8���Ћ���Qj�j��M�QP�΋RL�ҡ���H�A�U�R�Ћ���Q�J�E�P�у�_��^��]Å���   ��   vh����B�P�M�Q�ҡ���H�Aj j��U�h$SR����
����
�}�u�m�(S�M�Qj0j jj ���U��$R��������   ��|>��   v4����B�P�M�Q�ҡ���H�Aj j��U�h SR���m��땋���B�P�M�Q�ҡ���H�Aj j��U�hSR�Ѓ��M�Q�U�WR��������uPV�m������H�A�U�R�Ћ���Q�J�E�P�у�_��^��]���������������U��EHu�E�M�������   ]� �������������U��EHV����   �$���   ^]á��@�����uT�EP�7�����=�2  }�����^]Ëu��t�h4Sjmh��j��������t �����������tV���l����   ^]����    �   ^]ËM�UQR�V���������H^]�^]�ZU�����u.�ES������������t��蝑��V�׻�������    �   ^]Ã��^]�0�ɽн(��������h��Ph�f � ������������������U��h��jh�f ���������t
�@��t]�����]�������U��Vh��jh�f �����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R芐���E�NP�у�4�M��贐����^]ÍM觐�����^]��U��h��jh�f �\�������t
�@��t]��3�]��������U��h��jh�f �,�������t�x t�P]��3�]�����̋�3�� lS�H�H���������������̋A��t�x u3�ËQ����+����#�����������������U��E��x;A}
�I��]� 3�]� �U��E��x;A}�I�U���   ]� 3�]� ���������V��FW��u�~��N�<��u�< ��u_3�^á���H�F��  hpSj8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��S�]V��F;�~ ��x�F�M��^�   []� ^3�[]� }jW�F9FuK��u�~��N�<��u�< ��tA����B�V��  hpSj8��    QR�Ѓ���t�F�~�N�V��    �F9^|�_�F;Fu���������u����N�V�E���   F^[]� ��U��V��FW�};�~����y3�;Fu�m�����u_^]� �F;�~�N�T����H�;��F�M���F_�   ^]� ����U��E��x2�Q;�}+J�Q;�}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�C���3����_�F�F^�����A    ��������̋Q�B���x;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�A�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W��S�M���3����_�F�F^��������������U���SV�uW���^S�}�����3���F�F�O�N�W���V�E9G~|��I �O���F�U�9FuL��u�~��~��t���< ��tY����H���  hpSj8��    RP�у���t0�~�}���V��M����E�F@�E;G|�_^�   [��]� _^3�[��]� U��V�u��x'�A;�} �U��x;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��x,�Q;�}%��x!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|����Ѕ�x);�}%N�q;�}�A�t���B�0;Q|�_�   ^]� _3�^]� ������U����E�Qj�E��ARP�M��E��S�{�����]� �����U����Q�Ej�E��A�MRPQ�M��E��S������]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�lS��t!�A��t�B�A�Q�P�A    �A    �̋�� �S�@lS�HV3��q�q�P�r�r�lS�p�p�p�P�H^������V����S�r����F3��FlS;�t�N;�t�H�F�N�H�V�V�F�FlS;�t�N;�t�H�F�N�H�V�V^�U��U�E�V�2�0�
^]������������U����M� �S�H]� �����������U��E�UP�AR�Ѓ�]� ���������U��V��N3��lS;�t�F;�t�A�F�N�H�V�V�Et	V薱������^]� ������������U��V��W�~W��S�*���3����E��F�Ft	V�Q�����_��^]� ������U��V�������Et	V�)�������^]� ���������������U��Q�U�MSV�uW��y7��U��߃���   ����������U�A�Q����Q����Q��Q
����A����Q	����Q��Q����A����Q�������+�+�+�Ë���3�+�����3�+�+�����3�+�+ǋ���3�+�+��Ѓm���3�+�+�����3�+�+ǋ���3�+���+���
3�+���+���3���M�+����U�E�H��
wc�$����A
����Q	����A����Q����A����Q����A��Q����A����Q�����+�+�+�����3�+�����3�+�+����3�+�+�+�����3�+�����3�+���+���3�+�+ߋ�+���3�+�����
3�+�+���3�_^[��]Ë�1�(�������������������U��E�M;�}��]����������������U��E�@� �@����������������]��W  �����������̋���������������U��U���M��M�P�U�H�P]� U�조��Pl�E�I�RP�EP�EPQ�҃�]� ���������U��M�E���A�X���X]�������U����U�����Au���A�Z����Au�B�Y�A�����z��Y�A�Z����z�B�Y]� U��E�@� �@����������������]�U���8�E�M�� �A�`�A�M�`�� �A�`�A�M�`�� �]��A�`�]��A�`�]����������������������������������E����E������]��E����E��������]��E��������]��������������8V  �]��E����E������E������V  �E���P��]�U��E�M�� �A�`�A�M�`�� �A�`�A�`�������������������������������������������U  ��P]��������������U��E�H�P;�u'�I�M��R�P� �R�э@R��Q�^�����]�V�4R�U�I�ʍ4�VQ�H� �I��Q�@��Q�_�����^]����������U���h�U�J��RV�u�I�΍΍@�$ƍƍR�U��A�`�U��A���`�U��� �U��A�`�U��A�`�U������������]������������]������������������]������]����]��E����E������������T  ��P�]���W�qT  ��W�M��E����E������E������E����E�^�����E��������E����E������E�����������]�����U��A�M��%���]� �����������U��A�M��%   �]� ����������̋A$�������������U��E�M��V�uA������M�^]����������������U��E�M�US�W;�u;Pt�x;�u
;�u_3�[]�V;�u;Pt�p;�u;�u
^_�   []�;�u;Pt�@;�u;�u
^_�   []�;�u;�t;�u;�u
^_�   []�^_���[]��������U��E���T  �$�H��E��M��P�Q�P�Q�P�Q�P�Q�P�Q�P�M��P�Q�P �Q�P$�Q�P(�Q�@,�A]ËE�P�M��P�Q�P �Q�P$�Q�P(�Q�P,�Q�P0�M��P4�Q�P8�Q�P<�Q�P@�Q�@D�A]ËE�P0�M��P4�Q�P8�Q�P<�Q�P@�Q�PD�Q�PH�M��PL�Q�PP�Q�PT�Q�PX�Q�@\�A]Ã} �E�H0u�HH�UV�1�2�q�r�q�r�q�r�q�r�I�J��M��P�Q�P�Q�P�Q�P�Q�@^�A]ÍI ��F�������������U��E�H3�;H��]������������U��E��wM�$����E�M�]ËU�E�P]Ã} t�E�M�A�A]ËM�U�J]Ã} �E�Mt�A�A]Ë�������������U��E�M��]���U��E�M��]���U��E����   �$����M�E���Q�P�Q�P�Q�P�Q�I�P�H]ËM�E�Q��Q�P�Q �P�Q$�P�Q(�I,�P�H]ËM�E�Q0��Q4�P�Q8�P�Q<�P�Q@�ID�P�H]ËM�E�QH��QL�P�QP�P�QT�P�QX�I\�P�H]���E��P�X]�&�P�{���U��E�H3�;H�B]�����������U��M�E;u,�M�    �P3�;P�U�E�����
�    �   ]�;Hu"�M�U�E�   �    �    �   ]�;Hu+�M�U�   �   �H+H�U��Ƀ��
�   ]�;Hu"�E�M�U�    �   �    �   ]�3�]������U���S�]W���.����M���$���;�t_3�[��]�V3���~A��E�P�M�Qh���V���۶���M�U�R�E�Ph���V�Ŷ���M�;M�u�U�;U�uF;�|�^_�   [��]�^_3�[��]������������U���   �E��PSV�p�@W�u��u܉uȋu�E�E��E�EЉEԍE��VP�]��U��UĉU�M��M�M؉U������]��M�VQ�����E��U�VR�]��z����]��E�VP�m����E��M�QV�]�������]��U�RV������M��E�PV�]������]��M�QV�����M��E�P�	   ����|����M��@�`t������|����p�1`t�����}��p�1`t�����u��@�`t�����M�;�u���u	;�u	���t3���   ;�u���u	;�u	���t3���   ��t7����   �E����E���������������W����zq�����U�����{l�E��W�U؉�U܉P�U��P�U�P�E�Uȉ�ỦP�UЉP�UԉP�E �U$�    `���   ���{n��tj_^�   [��]�������Au��E�؋M���W�U��]���H�MĉP�U�H�E�M��U��H�M�P�U �H�E$�    �    @����Au�_^3�[��]�������U��U��VW�E�P�M�Q�MR3�W3�������tHS�U��M�G;�"�]���+ʍD�A��3�;P�Ã�C�Iu�U�E�P�M�Q�MRW�ȳ����u�[_��^��]������������U���W�E�P�M�Q�Mh���3�W葳����t/�E��M�G;�
��0@;�~��M�U�R�E�Ph���W�b�����u�_��]����������U���h��S�]�U�V�UЋu�U؋V�U�W�U�E��U�P�U�3��U�;V�U��M��U����U�Q�]��MPQS������<�C�����uVSW�H������U��H�����U��M�Q�N�U�R3�;N�M��RQP�����E���4;�uO;]�uJ�E��e��E��e��E��e��E��������������������������A��   �E��e��E��e��E��e��M;}�uo;�uk�E��e��E��e��E��e��E��������������������������Au7�E��e��E��e��E��e�����������������������z_^�   [��]���_^3�[��]��̋�3ɉ�H�H�H�H�H�H�H �H�H$���������������V��V�G����FP�>����NQ�5����VR�,����FP�#����NQ�����V R����3����F�F�F$^��U��E;A$|3�]� �QV�4��U��1W�2�q�|�+<��4��z�q �4��y�4v�4��r�q �4���q�r�q �4�q�r�q �|�+<��4��z�q���I��_�B�   ^]� �����̋�3ɉ�H�H�H�H�H�H��������U��E=   @w?t$��t=    up�E�@   �     �@   ]ËE�    �@   �@    ]�=   `t =   �u0�E�    �@   �@   ]ËE�@   �     �@   ]�����U��QSW��3�9_~a�]�V�W���E��O��������   ��4v��uVR�P���R�P���R�P� �����R�P�#  �E�C��;_|�^_[��]� ��������U���d��S�U�V�U���M�U��U��U��U��U��U��U��U��U��]��^��3ۉE�9^��   �]W��    �F�<�����QD�M��R,�E�P�����WQ�ҋE�N�U�R�V����   �R�P���R�P���R�P� �����R�P��"  ����QD�M��R0�E�PWQ�҃EC��0;^�t���_^[��]� �����������V�q3ҋƅ�~�I��tHB;�|�^���U��VW�}3�9w~S�]�G�������Q��詭��F;w|�[_^]���������������U��j h*  �a����������   �M�R|Q���ҋ�QU���F��]� ��������U���$  �MSV3�W�]��w\���u�}�M$�E��E �������  9]��  ����B���   h�W����h-  Q�҃������  ��~2ǅh�������3ɋא������8��x����x��h�����J�xu�3��}�9]��  ����Hl�I�U�R�U�E�P�BWP��3ۃ��]�9]��R  �����ݕ����������ݕ����Qݕ���ݕ���ݕ���ݕ���ݕ$���ݕ,���ݕ4���ݕ<���ݕD���ݝL����BD�U���U��@,QR�ЋM���U�6�����A3�;A�E���P�E����UԍU�RPQW�����U�������QR��T���P����3���,�}؉}����  ��I �}�����ݕt�����t���ݕ|���P�U��U��U��U��U��U��U��U��U��]̋QD�M���M��R,PQ�ҋE�<���l���Q��p���R�U����M�E�PQR�����]܍�t���P������SQ������ ܥT�����,�@ܥ\�������������W����AtF�E������U�3Ƀ}��E�   ����w#�$������F��F��u	�
��t�F�F�E�@�E�;E�������}� �]�uV�M�3��}�����wB�$����U���4�E��F�,��t�E��F�F��M��N���t�E��F�F��U��V�E��}�uC�]�;]������G�}�;}�s����]��M��~u�E�����+Ѝx�U܉M���I �U܋�ǃ8 }�C�x }�XC�x }�3�;O�X�ʅ�t�XC�x }�3�;O�X�ʅ�t�XC���M�u��E$�����Q���   �[�h�W��hi  P�ыU 3Ƀ��;�u$V赕���E P謕���M$��_^�����3�[��]ÉM$9M��   �M��	��    �u�]�3��S;S��3��x����   ����ݕt�����t���ݕ|���P�E��U��U��U��U��U��U��U��U��U��]̋QD�M$Q�J,P�э�t���R������VP�������U ��I�ʋ��P�Q�P�Q�P�Q�P�Q�@F���A;��g����E$�E�@�E$;E�3���_^�   [��]ÍI s�w�|���������������V��蘧���F�    ��^�������������    �I�R�����U��E�U	�IR�ܧ��]� ��������U��U�HX��S�V�u�Z3��@X�R�Z9^~[W3����N��9�����Au���B�Y����Au�A�Z�B�����z��Z�B�Y����z�A�ZC��;^|�_^[]�������U��E���$SV�uW�}����T�3�;T�������E�Ӄ�w/�$�8��U ��!�U �P��ҋU �Pu��ҋU t�P�P�E������������U�8���M��]�}��E�    �U�t�E$�����Bl�M�Q�@WR�ЍM�Q�U�R�U��M�QVPRWS�c+  �E��E����Ql�E�H�R��(WQ�ҋM�����y� �
�D��M��}�U�;���   �`��   ����   �����E�P�M�Q�U�RVS������F3҃�;F�E�@�u��    �����E��w/�$�H��U ��!�U �P��ҋU �Pu��ҋU t�P�P�E��t�E$�����Ql�E�H�RWQ�ҋu�]�M�Q�U�R�U��M�QVPRWS�S*  ������M$��$;��M  �E��U�E��E������<�����E��E�E�    �Ql�H�RWQ�ҍM�Q�U�R�U��M�QVPRWS��)  ����Hl�U�B�I��(WP�ыM�����y� �
�T��E��}�;}���   �`��   ����   �����U�R�E�P�MQVS�x����V3���;V�u����    �ЋE�@���E��w/�$�X��U ��!�U �P��ҋU �Pu��ҋU t�P�P�E��t�E$�����Ql�E�H�RWQ�ҋu�]�������M$��$_^[��]�,�3�;�G�_�f�n�z�����������������U��j�hzd�    P���   SVW��3�P�E�d�    ����3ۉE��]��E�@$�]��]�;���  �U�M�Q�MR�]ȉ]Љ]ԉ]܉]������E܋}�PW��������QHS�����   h�  V�Ћ���QHS�E苂�   h�  V�ЉEă� 3��ω}�;�~���U��tI@;�|�M�9]�~0�M�UȋE�+щE�
��D
�A�D
�A�D
�A���M�u�;�~6��E���X�M����A���A���O�����������X��X��X�u����؋���Q�J��|���P�ы���B�PSj���|���h�XQ�ҋE�P��,���Q�E��y�������������   �M�Px�E��ҍ�|���QP�����R�B��WP��<���P�E���A����������   P�B|���E��Ћ���Q�J��<���P�E��ы���B�P�����Q�E��ҡ���H�A��,���R�E��Ћ���Q�J��|���P�]��ы���B�P��d���Q�ҡ���H�ASj���d���h�XR�Ѓ�$Sh*  ���E�����������   �R|����d���P���ҋ��I����x�������H�A��d���R�]��Ћ���Q�J��L���P�ы���B�PSj���L���htXQ�҃�Sh*  ���E�莬����������   �R|��L���P���ҋ��|H����`�������H�A��L���R�]��Ћ���Q�J�E�P�ы���B�PSj��M�h`XQ�҃�Sh*  ���E�������������   �R|�E�P���ҋ�� H���E�����H�A�U�R�]��Ћ���Q�J�E�P�ы���B�PSj��M�hPXQ�҃�Sh*  ���E�虫����������   �R|�E�P���ҋ��G���E�����H�A�U�R�]��Ѓ�3�9]�~P�MԊ9�E�t��x���W�`����E�t��`���W�M����E�t	�M�W�=���;}�}	�M�W�/���G;}�|�������   �PSj���ҋMSSSV�����E�M@�E�;A$�����S��&���U�R�E������n������M�d�    Y_^[��]����������U��j�h�d�    P��SVW��3�P�E�d�    3�9]tX�u;��  ���?������  �};���   �EP�M�]�]��  W�Ή]�������E�;�u#�M��E������  3��M�d�    Y_^[��]�3�;�~=�M��8t*�A�u����u���A��u���A��u���E�B��;�|�3�;�~A�M�U���I �Y��< u�Y��< u��< u	�Y�< t
��U�E�F��;�|ˋMWP�!����M�Q�����U�R�E������؉������M�˝���   �M�d�    Y_^[��]�����U��j�hd�    P��   SVW��3�P�E�d�    ���}�3��w�7�w�w�w�w�w�w �w9u ��  9u$��  �m����E��]�u�;�t$��虜����~��莜��;E �E�P��讝����M IQ�M�V�Μ��9u,��   �}  �E    ~l�u�����F��;�t:�^;�t3�V;�t,;�t(;�t$��x ��x��x��x�]$;�};�}	9^};�|�E,�U�H�R�;����E@���E;E |��E,�8 ��  �M��؛���] �US�E��E�RP�����M���S��Q�Mĉu��  3�V�M��E��]��]��  �UR��P�M��E��]܉]��]��]��]�  ��t"�E�;�}�M�Q�M�����R��R��  ���]��E��PQ�M��E��]܉]��]��]��]��  ��t"�E�;�}�U�R�U�����Q��P�  ���]��E �M$���E�;�}��P�M�]�]��w  �u��E�9]���   9]���   �M�Q�E��a������]�]��E�;�~�U��E,P�U,�A������E�9]�~�M��U,R�M,�&������E�P�E������]��]�M�Q�E������U�R�]̉]��E� ������E�P�]ĉ]��E������
�����3��M�d�    Y_^[��]�( 9]��J���9]�u	9]��<���9]�u;��/���9]�u
9]�t� ���9]������M��  ������3�3��M��uԉ]܉]�蠰���E��w����E�M��U P�EQ�M$RPQ�E�����������   �UR�E��R������u�M��E��`����M��E���  �M��E���  �M��E���  �M��E��p  �M��E� �T  �E�P�E������������3��M�d�    Y_^[��]�( �}, �C  �M,�U�E Q�MR�U$PQR��#  ������   �E��EP蠘�����E    �M��E�誯���M��E��>  �M��E��B  �M��E��6  �M��E��  �M��E� �  �M�Q�E������>�����3��M�d�    Y_^[��]�( �U,�: ��   �EP�E��������M��E    �E������M��E��  �M��E��  �M��E��  �M��E��&  �M��E� �
  �M��E�����Q誗�����   �M�d�    Y_^[��]�( �U�E �MR�U$PQR�M�趮���E���������UR�a������} t#�M耗����~�E�u�P������uԋ]؃��} t#�M�W�����~�M�u�Q������uԋ]؃��U R�M��E     �	  �E P�M��E     ��  �}� �f  �F���}�E$;���  �����E��EE�����ɉH����HɉH�EċMԋ��������MP�M �@��M�E��M�Jl�U��AR�Ѓ���3���u�E �H;H��   �D��M��� ���   �������   �U����1��   ��W�Ũ����$��E�[��M�<��P�E Q�MVPQu)���������t�T��E�@�y   �D��U� �l��������u�T��E� �S�D��U���E̋��E$;]|;�|6�Mċ����M$�M̉��M$�U��Ủ��Uĉ��MċU���@�E$�� F��������EԃE@�E�;E$������}3�;}$��   �U���Eċ���E3ۋH;H�ÍK3ۉM��~[�����E��I �< }=�E#P�E�V�M�QP�E�M�QWPR���E# �����E�U؊M#��U��M�E�� FC���E;�|�G;}$�x����]��E܍U$�R�M��]��1  �E�P�M��%  �u�;u�������}��E��M܉�E��O$�M�3��G�E��O�_�G ����u��u�B���   h�W��hS  Q�u��u��u��u��u��u��҃��G;����������Q���   h�W����hT  P�у��G;�uq�M��E�������M��E��  �M��E��  �M��E��  �M��E��  �M��E� ��  �U�R�E�����苓����3��M�d�    Y_^[��]�( ����H���   �[�h�W��hU  R�Ѓ��G;����������B���   h�WhV  S�у��G;��3����u��u��u�3��E�	�E$9w$�  �O���w �����I+ʉM܍��p����O�U �MԋO�[�ыM ����+�}( �]�U؉M�}���  �E��E    �u;�u�}� D;��E~�E��MQP�M��D  ���c  �E�;�~�UR�U���+�Q��P�   ���M�u��U��F��E3��E    ��~?��U��M���t�M��I�M�
�M��A�M�M��Ȋ��@�;�|ƋM�E܅���  �U �҉U ���E�G3�;G��3��A�E����   ���U����M ���Eċ�@��U��l���RVP�����݅l����UԋM �����݅t����\��Eċ���E���U�@�ʋU؍[�ʋ��P�Q�P�Q�P�Q�P�Q�@F�A;u�g����}u�O�O�E ���M�0�����   �U܅���   �} ��A��E �U3ۍ�    �3�;P����;���   �E �t���Mċ�@��U��l���RSP������ �@������Eԃ���X�Mċ�M�����@�E�ЋU؍v�ʋ��P�Q�P�Q�P�Q�P�Q�@�U�A�M�Ί�M�$��E C�Q��������M�E �7����E$�U�@�E$;B$}�������M��E���  �����}, �u�tf3�9^$~_�N ����3�;A}�V �T��N�tG@;�|��}.�F�<�;|���}�Mċ��M,�	�IP�	����VG;|�|�C;^$|��M��}�O�F$�V���Y���  �������E�����E$�����E ��    �E 3ҋH;H�ʅ�tr�U�N �
�V�I��QP�!  ���}, t��t�Uċ��E,�H�R�o�����E ��M$��P�Q�P�Q�@�A�Mċ��V%�������   �Eċ��UR�EP��t���R�U荅\���P�F R�U��V�@��PQ�M��<����M PQ� ����� ���@�}, t��t�Uċ��E,�H�R�Ɏ����M$��\������`����T��d�����P��h����P�Eċ��U3�%���3V�����x�������M$��t������|����P�U��H�M�P�Eċ�3�K%���3��N���V�E;<u�m��   )E )E$KO�]����M��E��q  �M��E�赤���M�Q�E��Xz��3����M��u�u��E��A  �M��E��5  �U�R�E��(z�����Mĉu��u��E� �  �E��E�����P�������U��Q���SV�uW���HH���   h�  V�ҋء���HH���   h�  V�҉E����HH��p  j h�  V�҉E�����HH��p  j h�  V�ҋM �U��(Q�MR�USQ�MR�UQ�MR�U�QRP������_^[��]� �����������U��j�h1d�    P��SVW��3�P�E�d�    �M���HH�]���   h�  S�҃�3�P�M�u�u��
  �M�u���;���E����HH���   h�  S�҃���~H3��	��$    ���E����QD�J,�P�EVP�ы���BH���   h�  SF��`�у�;�|ŋU �E�MR�UP�EQ�M�RPQ�M�S�d����U�R���E������Rx�����ƋM�d�    Y_^[��]� ���������U��E��PVW;�tB�x;�t;�@;�t4;�t0;�t,��x(��x$��x ��x�u;�};�};�};�}	_�   ^]�_3�^]��������U��E�MPQ�������W������z�   ]�3�]������U��E=   @��   ty��t9=    ��   �E�M���A�M�X��X�A�M�X ��X0�A�X8]ËE�M���A�M�X��X�A�M�X ��X0�A�M�X8��XH�A�XP]ËE� �M�YH�@�YP]�=   `t=   �u?�E� �M�Y0�@�Y8]ËE�M���A�M�X��X�A�M�X ��XH�A�XP]���U��E�MP�E�P��Q�M�R�P���R�P� �����R�P�������]���U���E����X]� ���������������U���E����E�X]� ������������V���H������^���V��V�G������    ^������������̋�������������̋��������������U��E]� ���̃9 u�y t�   Ãy ~�3�������̃9 u�y t�   Ãy ~�3��������U��E��]� ̃9 u�y t�   Ãy ~�3�������̋�    �A    Ë�3ɉ�H�H���̃9 u�y ~�   �3��������������U��E�@��]� ��������������U��E]� ����U���M��]� �U��E��]� ̋3҉�Q�Q����U���M��]� �U��E�@��]� ��������������U��V�uV�t�����    ^]� �����U��V�uV�ct�����    ^]� �����U��V�uV�Ct�����    ^]� �����U��V�uV�#t�����    ^]� �����U�조��H�U����  hOh5  P�у�]� ������U�조��H�U����  hO��h5  P�у�]� ��U�조��H�U����  hO��h5  P�у�]� ���U�조��H�U����   h�N��j!P�у�]� �����U��V�u��MQ�E�;s�����    ^]� �������������U���E� O�  ]� �����������U�조��H�U����  hO�@��h5  P�у�]� U��E��t	�M��]�3�]��������������������������U��M�E���A�X]�������������HX��Y�@X�Q�Y��������̃9 u�y t�   Ãy ~�y u�y t�   Ãy ~�3����������������V�qV�F������    ^������������U��E]� ����U���M��]� �U��E��]� �U���M��]� ̋3҉�Q�Q����U��E�@��]� ��������������V��V�q�����    �F    ^������V��V�gq�����    �F    ^������V��V�Gq�����    �F    ^������V��V�'q�����    �F    ^������U��V�uW��9wu_�   ^]� ����H���  ShOh5  V�ҋ؃���t=��~9�G��;�|�ȋ��t��tQPS��  ���G;�~��+�Q�j P�W  ��W�p������w��t��u	[_3�^]� [_�   ^]� ���������U��V�uW��9wu_�   ^]� ����H���  ShO��    h5  R�Ћ؃���tG��~C�G;�}�ƍ�    ���t��tQPS�4  ���G;�~��+���Q��j R�  ��W��o������w��t��u	[_3�^]� [_�   ^]� ��������U��V�uW��9wu_�   ^]� ����H���  ShO����h5  R�Ћ؃���tD��~@�G;�}�Ƌ����t��tPQS�z  ���G;�~��+���Q���j P��  ��W�o������w��t��u	[_3�^]� [_�   ^]� �������������U��V�uW��9wu_�   ^]� ����H���  ShO�v��h5  R�Ћ؃���tM��~I�G;�}�Ƌ�@����t��tPQS�  ���O;�~��+��@���IR���j P�  ��W�Hn������w��t��u	[_3�^]� [_�   ^]� ���U��E�U����;�sV�uW��t�>�9��;�r�_^]�����������������������U��E�U����;�s V�uW+���$    ��t�<�9��;�r�_^]�������������U���ES�YV�4�W�}���<��Y�������4�_^[]� ���������������U���M��]� �U��A�M��]� U��EV��P�    �F    ������^]� �������������V��V�m�����    �F    ^������U��EV��P�    �F    �t�����^]� �������������V��V�l�����    �F    ^������U��EV��P�    �F    �������^]� �������������V��V�gl�����    �F    ^������U��EV��P�    �F    �T�����^]� �������������V��V�l�����    �F    ^������U��S�]�V��;Fu^�[]� ����Q���   Wh�N��j!P�ы�����t?��E�RQW��������~ ~��EP�U�k�����    �>�_�N^�[]� _^2�[]� ��������U��QV��~ ~��M�Q�E��Uk�����    �    �F    �F    ^��]����U��QV��FW�~;F}�����t�U�
���P�_^��]� @�E��E�� O�l  �E��E�PW���������u_���^��]� ������t�M����H�_^��]� �������������U��j�hcd�    P��SVW��3�P�E�d�    ���}�3���G�E��G�G�M�E��}��P��������uV�O������? u� t�   � ��   � u� t�x   � ~r3���~�O������@;�|�M�U�R�E�Ph���3�V�E    �>~����t:�E��E;E�����W�4�@F;E�~�U�E�P�M�Q�Mh���R�~����uƋǋM�d�    Y_^[��]� ����������U��j�h�d�    PQVW��3�P�E�d�    ��u��~W�E�    �Fi��V�    �G    �E������,i�����    �F    �M�d�    Y_^��]������������U��QV��~ ~��M�Q�E���h�����    �    �F    �F    ^��]����U��EVP�������> u�~ ~�   3Ʉ���^��]� 3�3Ʉ���^��]� ���U��SV�uW���G;�u� L�} u;�~?;��E~�G�MQP���H�����u_^[]� �G;�~�UR���+�Q��P�������w_^�[]� ���U��SVW�}���    �F    �F    �}�E��~�F�MQP���������t!�F;�~�UR���+�Q��P�������~_��^[]� ����������U��} ���ЋER�UPR������]� ��������������U��M�U$�ESV�u ������M�������E������UW�}9zt9t9Hu�    �T9zt9Ht9Hu�   �=9zt�X�x;�t;�t;�u�   ��}9zt9Ht9u�   ��> |��L��E$�����E�_^[]����������U��E�M S�]V�uW�}� ���������3ҋ�����ǅ�x;Mt90t9pt9pt9ptB��|�_^[]ËE_��M ^�[]��������������U����E��U�j �M��M�jQ�E��M�������]�������U��E�VW��xE�p��x>�x��x7�@��x0�M;�});�}%;�}!;�};�t;�t;�t;�t;�t	_�   ^]�_3�^]��������U����E�Mj �U�jR�E��M������3҃��u��]���̃9 u�y t�   Ãy ~�3�������̋A������������̃9 u�y t�   Ãy ~�3��������U��E�	����]� ��������������U���M��]� �U��V�uV��d�����    ^]� �����U��V�uV��d�����    ^]� �����U�조��H�U����  ��hO��h5  P�у�]� ���������������U�조��H�U����  hO��h5  P�у�]� ��U��E�	����]� ��������������U���M��]� �V��V�d�����    �F    ^������V��V��c�����    �F    ^������U��V�uW��9wu_�   ^]� ����H���  S��hO��h5  R�Ћ؃���tM��~I�G;�}�Ƌ������t��tPQS�  ���O;�~��+�����R����j Q�  ��W�Gc������w��t��u	[_3�^]� [_�   ^]� ��U��V�uW��9wu_�   ^]� ����H���  ShO��    h5  R�Ћ؃���tG��~C�G;�}�ƍ�    ���t��tQPS��  ���G;�~��+���Q��j R�V  ��W�b������w��t��u	[_3�^]� [_�   ^]� ��������U��EV��P�    �F    �d�����^]� �������������V��V�'b�����    �F    ^������U��EV��P�    �F    �������^]� �������������V��V��a�����    �F    ^������U��j�h�d�    P��,SVW��3�P�E�d�    �}3�;�t����t������u��    P�MЉ]Љ]�������    Q�M؉]��]؉]��2����E�9]�u?9]�t?�M�Q�E� �7a���U�R�E������]؉]��!a����3��M�d�    Y_^[��]�9]�~�9]�u9]�t�9]�~�3��]�E�;�t%�UR���-v���E�;�u�E�P�E� ��`���M�Q�3ɉM9]��  �u���u�;�t
�< �d  �N�;�|;�~�;�|4�^���x-���x'�E;�} ;�};�};�};�t;�t;�t;�t;�u�U�MjR������E��3����M��E���u�F�;��   �D��A���L���;�|C���؋u�j �M�jQ�}ȉ]��0���3����M؃��<� t%�u܋�98u9Xt�F�;�}B����3҃<� uދ4���u0�EЋu�Ɖ��U�   M���u��P�@�����H�8�X�?�~u�E�F�F   �*�N�}jQ�������VjR�������EjP�������M��u�A�M��������E�M3�A���M�u�;M�{���;�t�M�Q�_�����U�R�E� �
_���E�P�]؉]��E�������^�����   �M�d�    Y_^[��]ø�3�����*��?*��x*���)��� �j3�$��)�(�_)�,��(Ë�U��M������]Ë�U�������} t��  ��]������������̋T$�L$��ti3��D$��u���   r�=�� t��  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u�  ��   u������r)��$�@�Ǻ   ��r����$�T�$�P��$���d��#ъ��F�G�F���G������r���$�@�I #ъ��F���G������r���$�@�#ъ���������r���$�@�I 7$���D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�@��PXdx�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$���I �Ǻ   ��r��+��$���$����<�F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ���������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U���uQ�^  YY]� ��Q��X��  YË�U��V��������EtV�b]��Y��^]� ��U���uQ�  YY]� ��Q��  YË�U��E��	Q��	P��  ��Y�Y@]� ��U��E��	Q��	P��  ��Y�Y��]� ��U��E��	Q��	P�  YY3Ʌ�����]� �AË�� �X� ��� ��̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$���58������t��j��  jj �~  ���C  ��U��V�58�����u������8���^]��58�����;�u���   jh���2  �E��uz��1  ��u3��8  �$  ��u��1  ���X1  �������0  �����*  ��y�J!  ����/  ��x �N-  ��xj �l(  Y��u�����   ��,  ��3�;�u[9=��~�����}�9=��u�4*  9}u�,  ��   �51  �E������   �   3�9}u�=4��t�   ��j��uY�\   h  j��%  YY��;�����V�54��5l�����Ѕ�tWV�   YY�����N��V�C  Y�������uW�#  Y3�@��0  � jhУ�0  ����]3�@�E��u9����   �e� ;�t��u.��X��tWVS�ЉE�}� ��   WVS�C����E����   WVS�����E��u$��u WPS�Ԝ��Wj S������X��tWj S�Ѕ�t��u&WVS�������u!E�}� t��X��tWVS�ЉE��E������E���E��	PQ�b3  YYËe��E�����3��0  Ë�U��}u�]3  �u�M�U�����Y]� ��U��QSV�5��W�5�����5���؉]��֋�;���   ��+��G��ruS�3  �؍GY;�sH�   ;�s���;�rP�u��9$  YY��u�C;�r>P�u��#$  YY��t/��P�4��������u�=���׉��V�ף���E�3�_^[�Ë�Vjj �#  YY��V�����������ujX^Ã& 3�^�jh��.  �$  �e� �u�����Y�E��E������	   �E���.  ��g$  Ë�U���u���������YH]Ë�U��=�� u�_  j�  h�   �
$  YY�E��u@Pj �5�����]Ë�U��S�]���woVW�=�� u�  j�_  h�   ��#  YY��t���3�@Pj �5���������u&j^9��tS�3  Y��u���s2  �0�l2  �0��_^�S�3  Y�X2  �    3�[]Ë�U��} t-�uj �5�������uV�'2  �����P��1  Y�^]����̃��$��6  �   ��ÍT$�6  R��<$�D$tQf�<$t�P6  �   �u���=�� ��6  �   � ���6  �  �u,��� u%�|$ u���%6  �"��� u�|$ u�%   �t����-�c�   �=�� �f6  �   � ��o5  ZË�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$��XY�$��XY�$����U��QQSVWd�5    �u��E�$j �u�u��u�� �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u��G  �� �E�_^[�E���]�U���SVW��E�3�PPP�u��u�u�u�u�G  �� �E�_^[�E���]�U���SVW��E�3�PPP�u��u�u�u�u�WG  �� �E�_^[�E���]Ë�U��E�p�p(j �p��6  ��]� ��U��V��u�N3������j V�v�vj �u�v�u��F  �� ^]Ë�U���8S�}#  u��%�M�3�@�   �e� �E�&���M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��o  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M������E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u��E  �� �E�x$ u�u�u�q���j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����+���u�F  �MN��k�E�9H};H~���u	�M�]�u�} }̋EF�0�E�;_w;�v�KF  ��k�E�_^[�Ë�U��EV�u��  ���   �F��  ���   ��^]Ë�U����  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�  �u;��   u�  �N���   ^]��  ���   �	�H;�t���x u�^]�E  �N�H�ҋ�U������e� �M�3��M�E��E�E�E@�E�%�M��E�d�    �E�E�d�    �uQ�u�E  �ȋE�d�    ���Ë�U��]��E  ��U��EV���F ��uc��  �F�Hl��Hh�N�;��t�P��Hpu�O  ��F;X�t�F�P��Hpu�G  �F�F�@pu�Hp�F�
���@�F��^]� �y t�A�`p�Ë�Ë�U��} t�u�u�u�u�u�Q  ]Ë�U���V�u�M��3����u�P��X  ��e�F�P�dS  ��Yu��P��X  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�X  �M��E��M��H��EP�Y  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�]  @PV�V�Z  ��^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M����}���3�;�u"�?*  j^�0�O  �}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�*  j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]h�XSV�<]  ����ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F���_t�90uj�APQ�X  ���}� t�E��`p�3������3�PPPPP��M  ̋�U���,��3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0�E^  ����u��(  ��N  ���m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q�\  ����t� ��u�E�j P�u��V�u��������M�_^3�[�U����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �'���9}}�}�u;�u#��'  j^�0�7M  �}� t�E�`p����  9}v؋E��� 9Ew	�'  j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V�@  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �]  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� ��\  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�������u�E�8 u���} �4����$�p���W�T\  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP�)[  0�F�U�����;�u��|��drj jdRP�[  0��U�F����;�u��|��
rj j
RP��Z  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U��j �u�u�u�u�u�o�����]Ë�U���SVW�u���w�ٍM�N������u#�\$  j^�0�I  �}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^��V  @PVS�xS  �0�������} ~QV�^��V  @PVS�TS  �E����   � � ������y&�߀} u9}|�}�}�������Wj0S��������}� t�E��`p�3�_^[�Ë�U���,��3ŉE��EVW�}j^V�M�Q�M�Q�p�0��X  ����u�D#  �0�H  ���lS�]��u�,#  �0�H  ���S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P�W  ����t� ��u�E�j VS���N�����[�M�_3�^������Ë�U��j �u�u�u�u�'�����]Ë�U���,��3ŉE��EV�uWj_W�M�Q�M�Q�p�0��W  ����u�f"  �8��G  ���   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW�:V  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u�b�������u�E�jP�u���u�u�f�����[�M�_3�^������Ë�U��j �u�u�u�u�u�������]Ë�U��E��et_��EtZ��fu�u �u�u�u�u�������]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u������u �u�u�u�u�u������]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3��������������(r�_^Ë�Vh   h   3�V��W  ����t
VVVVV�E  ^�f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U���j
������3��W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����jh��  j��W  Y�e� �u�N��t/�����E��t9u,�H�JP�B���Y�v�9���Y�f �E������
   ��  Ë���j�}V  Y�jh0��  �}3�9_��   h (  h�"h"S�G	PS�F�  ���E�;�u3��   P�Q  Y���N�E�<0 u�0;�w�Nj�W  Y�]�9_uVj����Y�؅�tH��V�����Y�G��t0�u�VP�{Q  ��3�;�u�G��E�H�K�X�QQQQQ�B  S�N���Y�u��E���Y�E������   �G�  Ë}j�U  Y�jhP��  j�gV  Y�e� �u�N��t/�����E��t9u,�H�JP�����Y�v�����Y�f �E������
   �  Ë���j�U  YË�U��f�} u�E (  �uh�"h"�u�u�u��  ��]�jhp��  3ۋu9^��   j�U  Y�]�9^��   h (  S��	VS���������}�;�uj��E�Ph�脯  ��3��   W�TO  Y���u���N�u���t�>�8 u�  ��j�^���Y��;�tJ�^S�N���Y����t3�u�SV��O  ��3�;�u�E�p�7�E�H�O�x�QQQQQ��@  W����Y�u�����Y�u�E������   �F�T  Ëuj��S  Y�jh����  j�T  Y�e� �E�p��t�~�6�H���V�B���YY�����E������   ��  �j�S  Y���������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�����&�  ��tj�z�  Y�0�tjh  @j�G>  ��j�  ̋�U��M�0��U#U��#�ʉ0�]Ë�U��3��M;�Xat
@��r�3�]Ë�\a]Ë�U����  ��3ŉE�SV�uWV������3�Y�����;��l  j褶  Y���  j蓶  Y��u�= ���   ���   �6  h�bh  ��W���  ������   h  �B�VSf�J������  ��uhdbSV�ŵ  ����t3�PPPPP�>  V葵  @Y��<v*V脵  �E����+�j��h\b+�SP蚴  ����u�hTb�  VW��  ����u������VW���  ����u�h  hbW�v�  ���^SSSSS�y���j������;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]��K  YP�����PV����M�_^3�[�������j�)�  Y��tj��  Y��u�= �uh�   �%���h�   ����YYË�U���   ��3ŉE��}�ESVW�}��x�����   ��t��� h�   ��|�����Q�u�uP軶  ������ub�����zuxVV�u�u��x���蔶  ����p�����tXFVP��  ��YY��tH��p�����t���S�u�u��x����Y�  ������tjV�  �3�YY;�u!9�t���tS�N���Y����M�_^3�[�����ÍN�QSVP�L�  ����u9�t���tS����Y3���WWWWW�M<  �}uH�5��3�PP�u��u�֋؅�tjS�'  YY���tSP�u�u�օ�u��7������' Y�p����} �f�����x��� j��x���P�E    P�u������<�����x�����c�����U��E�8�]Ë�U���(  �H��D��@��<��58��=4�f�`�f�T�f�0�f�,�f�%(�f�-$���X��E �L��E�P��E�\����������  �P��L��@�	 ��D�   �����������������������j輴  Yj ���h�b����=�� uj蘴  Yh	 ����P�����j �������� ��U���u�58�� ���]� �4�Ë�V�58�� �����u�5h������V�58�����^Ë�U���u�u�5l������]� �4����tP�5p�����Ѓ4���8����tP���8���L  jh���)  h�b���u�F\@c�f 3�G�~�~pƆ�   CƆK  C�Fh0�j�M  Y�e� �vh���E������>   j�M  Y�}��E�Fl��u����Fl�vl�4  Y�E������   ��  �3�G�uj�dL  Y�j�[L  YË�VW����54��������Ћ���uNh  j�  ��YY��t:V�54��5l�����Ѕ�tj V�����YY����N���	V����Y3�W��_��^Ë�V��������uj��  Y��^�jhؤ��  �u����   �F$��tP�<���Y�F,��tP�.���Y�F4��tP� ���Y�F<��tP����Y�F@��tP����Y�FD��tP�����Y�FH��tP�����Y�F\=@ctP�����Yj�&L  Y�e� �~h��tW����u��0�tW����Y�E������W   j��K  Y�E�   �~l��t#W�3  Y;=��t����t�? uW�*4  Y�E������   V�R���Y�  � �uj�J  YËuj�J  YË�U��=4��tK�} u'V�58��5 ��օ�t�54��58����ЉE^j �54��5l�������u�x����8����t	j P��]��%���%���Wh�b������u	����3�_�V�5 �hcW��h cW�d���h�bW�h���h�bW�l��փ=d� �5��p�t�=h� t�=l� t��u$� ��h����d�T?�5l��p�����8������   �5h�P�օ���   �q  �5d��5�����5h��d����5l��h����5p��l��֣p��rH  ��tc�=��hRA�5d����У4����tDh  j��   ��YY��t0V�54��5l����Ѕ�tj V����YY����N��3�@��]���3�^_Ë�U��V�uV�$����  ;5t�v�����^]Ë�U��M�t��t�]Ë�U��VW3��u�\�����Y��u'9t�vV�$����  ;t�v��������uʋ�_^]Ë�U��VW3�j �u�u�ʮ  ������u'9t�vV�$����  ;t�v��������uË�_^]Ë�U��VW3��u�u��  ��YY��u,9Et'9t�vV�$����  ;t�v��������u���_^]Ë�U��VW3��u�u�u�^�  ������u,9Et'9t�vV�$����  ;t�v��������u���_^]Ë�U��h(c����thcP� ���t�u��]Ë�U���u�����Y�u�(��j��G  Y�j��F  YË�V������V�  V�;2  V�����V��  V��  V�3'  ��^Ë�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��M��u�C  �    �3  jX]á����t�3�]Ë�U��M��u�  �    �i3  jX]á����t�3�]Ë�U��=�X th�X��  Y��t
�u��XY�����h$EhC�A���YY��uTVWh�O�p���� @�BY��;�s���t�Ѓ�;�r�=�� _^th��胯  Y��tj jj ���3�]�j h ��  j�TF  Y�e� 3�@9����   ����E����} ��   �5���5���֋؉]Ѕ�th�5���֋��}ԉ]܉}؃��}�;�rK�2���9t�;�r>�7�֋���������5���֋��5����9]�u9E�t�]܉]ЉE؋��}ԋ]���E�(F�}�4Is�E� ��t�ЃE����E�8J�}�<Ks�E�� ��t�ЃE����E������    �} u)���   j�TD  Y�u�@����} tj�>D  Y��  Ë�U��j j �u������]Ë�U��j j�u������]�jj j �������jjj �z�����Ë�U�������u�d���Yh�   ����̋�U���LV�E�P�8�j@j ^V����YY3�;�u����  ��   ����5d�;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5����@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9d�}k���j@j �����YY��tQ�d� ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9d�|���d�3���~r�E�� ���t\���tW�M��	��tM��uP�4���t=����������4����E�� ��E�� �Fh�  �FP�0�����   �F�E�G�E�;�|�3ۋ���5������t���t�N��q�F���uj�X�
�C�������P��������tB��t>W�4���t3%�   �>��u�N@�	��u�Nh�  �FP�0���t,�F�
�N@�����C���h����5d��,�3�_[^�Ã������VW������t6��   ;�s!�p�~� tV�<����@   �N�;�r��7������' Y������|�_^Ã=�� u�A)  V�5��W3���u����   <=tGV��;  Y�t���u�jGW�������YY�=����tˋ5��S�3V�;  �>=Y�Xt"jS����YY���t?VSP�P<  ����uG���> u��5���3����%�� �' ���   3�Y[_^��5�������%�� �����3�PPPPP�7-  ̋�U��E���]Ë�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF豬  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�̫  Y��t��M�E�F��M��E��詫  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9��u�&  h  ���VS����@�����5��;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H�|��5��3�����_^[�Ë�U���SV�L���3�;�u3��wf93t��f90u���f90u�W�=H�VVV+�V��@PSVV�E��׉E�;�t8P�8���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u�����Y�u�S�D��E��	S�D�3�_^[�Ë�V�ԝ�ԞW��;�s���t�Ѓ�;�r�_^Ë�V�ܟ�ܠW��;�s���t�Ѓ�;�r�_^�j h   j �P�3Ʌ����������5���T��%�� á������h�Pd�5    �D$�l$�l$+�SVW��1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋���t�O�30�e����O�G�30�U��������������̋�U���S�]V�s35�W��E� �E�   �{���t�N�38�����N�F�38� ����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t��褗  �E���x@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�}����E�_^[��]��E�    �ɋM�9csm�u)�=Td t hTd�C�  ����t�UjR�Td���M�U�D�  �E9Xth�W�Ӌ��F�  �E�M��H����t�N�38������N�V�3:������E��H���ږ  �����9S�O���h�W����  ������V9t�����   ;�r���   ^;�s9t3�Ë�U��V�/��������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U������e� �e� SW�N�@��  ��;�t��t	�У���eV�E�P�d��u�3u��`�3����3��\�3��E�P�X��E�3E�3�;�u�O�@����u��G  ����5��։5��^_[�Ë�U��} u�e   �    �%  ���]��uj �5���h�]Ë�U��E3�;̀�tA��-r�H��wjX]Ë̈́�]�D���jY;��#���]�������u��Ã��������u��Ã�Ë�U��V������MQ�����Y�������0^]Ë�U���m�����ujX]������M�3�]Ë�U��V�u��u
��$  jX��z���� �3�^]Ë�U���'�����ujX]��l����M�3�]Ë�U��V�u��u
�$  jX��G���� �3�^]Ë�U��E���]Ë�U��Vj�8  Y�5������u�����j����7  Y��^]�j �����Y��5�����Ë�U���5�������t�u��Y��t3�@]�3�]Ë�U��� �e� Wj3�Y�}��9Eu�����    ��#  ����x�MV�u��t��u�b����    �#  ����S�����E�;�w�M��u�E��u�E�B   �u�u�P�u���  ������t�M�x�E��  ��E�Pj 荣  YY��^_�Ë�U���uj �u�u�u�<�����]���������������̀zuf��\���������?�f�?f��^���٭^�����c�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����c�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����c���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�c��p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR誯  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��d�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��<d�����������,d�����   s��Ld��4d�����������$d�����   v��Dd떋�U��V�EP���ů  �\d��^]� �\d�	�  ��U��V���\d���  �EtV���Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR�7���YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =RCC�t=MOC�t=csm�u*�w������    �G  �f������    ~�X������   3�]�jh ��J����}�]��   �s��s�u��"������   �e� ;utb���~;w|�,  �ƋO�4��u��E�   �|� t�sh  S�O�t��N  �e� ��u��+���YËe�e� �}�]�u��u���E������   ;ut��  �s�����Ë]�u��������    ~�y������   Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�<���3�A��  ���3��jhH��)����M��t*�9csm�u"�A��t�@��t�e� P�q�����E������8����3�8E��Ëe��  ̋�U��M�V�uƃy |�Q�I�42���^]�����3�9��   ��Ë�U��EVW�}��tq�0��tk�>csm�u/�~u)�F= �t=!�t="�u�~ u�V������   �vW�1���YY�@������   �G�2������   �G�$������   ��O��O��������   �������    _^}��������    3�@]Ë�U��E��tA� �8csm�u7�xu1�H�� �t��!�t��"�u�x u�������   3�@]�3�]Ë�U��V�u�~��(  SWV�����} Y�csm� ���   �b������   98uu�S������   �xud�B������   9Xt(�2������   �x!�t�������   �x"�u,�
������   �p����Y��tj��������   ����YY��������   98uZ��������   �xuI�������   9Xt(�������   �x!�t�������   �x"�u�} t�������   �u����N���   �g����N_���   [^]�jX�jhh��Q����e� �M�U��u�����YËe��E������q����jh�������e� �u�UY��u��e���YËe��E������>����jh��������e� �u�U��u��3���YËe��E����������jhȥ�����e� �u�u�u�u�U��u������YËe��E����������Ë�U��3���;�u
�  �G  �E��E�9~OS�E�V�E�@�@��p� �M�q�P�GE�P�;�������u
K�������E��E�E�E�;|�^[�E���j��跫  ��������    t�  �e� ��  �M���  ������Mj j ���   �R�  ̋�SW3�3�9~�F�Lh�������uG��;>|�2�_[ð����U��V�uW��u�  �6��u�  �>csm�u�~u�F= �t=!�t="�t�q  �F�@�8�p�!��@�M��P����P����YY��tO�����3�_^]�3�@��j,h@������ً}�u�]�e� �G��E��v�E�P�����YY�E���������   �E���������   �E��������   �����M���   �e� 3�@�E�E��u�uS�uW�������E�e� �o�E�����Ëe��k�����   �u�}�~�   �O��O�^�e� �E�;Fsk��T;�~A;L;�F�L�QVj W��������e� �e� �u�E������E    �   �E��?�����E�맋}�u�E܉G��u�����Y������Mԉ��   ������MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v����Y��t�uV�F���YY�jhh��l���3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w��  YY����   SV��  YY����   �G��M��QP����YY���   �}�E�p�tH裩  YY����   SV褩  YY����   �w�E�pV��  �����   ���t|��W�9Wu8�V�  YY��taSV�[�  YY��tT�w��W�E�p����YYPV�  ���9��  YY��t)SV�#�  YY��t�w�'�  Y��t�j X��@�E���9  �E������E��3�@Ëe���  3��?����jh��������E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w�����YYP�vS�E�����FP�w����YYP�vS�$����E����������3�@Ëe��<  ̋�U��E����u��S�]V�0W�}��t� u!�=MOC���   =RCC���   ��@��   �>csm���   �~��   �F= �t=!�t="���   �~ u��������    ��   ��������   �F�@��   ��}�8�]��X���v�EP�E�P��������u
O������_�������   �} t]�u�E�P�uV�u������H=csm�u6�~u0�F= �t=!�t="�u�~ u�1������    u3���������   3�@_^[�Ë�U��} t�uSV�u�������}  �uuV��u 蛼���7�u�uV�����Gh   �u@�u�F�u�KV�u������(��tVP����]Ë�U���V�u�>  ���   W�������    tG�w������   ����9t3�=MOC�t*=RCC�t#�u$�u �u�u�u�uV�A���������   �}� u�O  �u�E�P�E�PV�u W艾���M���;M�sg���E�S�x�;7|G;p�B���H�Q��t�z u-�Y��@u%�u$�u�u j �u�u�u�u�����u�E����E��M����E�;M�r�[_^�Ë�U���4�MS�]�CVW�E� =�   �I��I�M����|;�|�  �u�csm�9>��  �~� ��)  �F;�t=!�t="��  �~ �  �������    ��  �
������   �u��������   jV�E�Ĥ  YY��u�  9>u&�~u �F;�t=!�t="�u�~ u��  �������    ��   �������   �����u3����   ����Y��u\3�9~�G�Lh��Ĳ����uF��;7|��3  j�u� ���YY�EP�M��Edd�   h���E�P�E�\d谣  �u�csm�9>��  �~��  �F;�t=!�t="���  �}� ��   �E�P�E�P�u��u W�F����M���;M���   �x�}�M��G��E�9��   ;O���   ��E�G��E��~r�F�@�X� �E��~#�v�P�u�E��r�������u�M��9E���M�E��}� ��.�u$�}��u �]��u��E��u�u�uV�u�����u�}���E��E����}�;E��P����}�} t
jV�����YY�}� ��   �%���=!���   �����   V�G���Y����   ���������������   �����}$ �M���   Vu�u��u$�C����uj�V�u�u�+������v�a����]�{ v&�} ������u$�u �u�S�u�u�uV������ �:������    t�T  _^[�Ë�U��V�u��詟  �\d��^]� ��U��SVW�������   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�M������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������ 3�@_^[]�jh��� ��������@x��t�e� ���3�@Ëe��E�����������9����������@|��t������jh�������5�������t�e� ���3�@Ëe��E������}����hm��������������U���SQ�E���E��EU�u�M�m�艡  VW��_^��]�MU���   u�   Q�g�  ]Y[�� ����U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�ݩ��3��ȋ��~�~�~����~����0����F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  ��3ŉE�SW������P�v�l��   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�������C����u�j �v�������vPW������Pjj �V�  3�S�v������WPW������PW�vS�	�  ��DS�v������WPW������Ph   �vS��  ��$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�˭����jh8��������������P��Gpt�l t�wh��uj ����Y��������j�x  Y�e� �wh�u�;5X�t6��tV����u��0�tV����Y�X��Gh�5X��u�V���E������   뎋u�j�&  YË�U���S3�S�M��*���������u���   �t�8]�tE�M��ap��<���u���   �p��ۃ��u�E��@���   ��8]�t�E��`p���[�Ë�U��� ��3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�`���   �E��0=�   r����  �t  ����  �h  ��P�x����V  �E�PW�l����7  h  �CVP�=���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP������M��k�0�u���p��u��+�F��t)�>����E���\�D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C��d�Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����95���T�������M�_^3�[�ª���Ë�U���j �M��Ǵ���E�x t�}� �@t�M��ap��À}� t�E��`p�3���jhX������M���������}������_h�u�3����E;C�W  h   �����Y�؅��F  ��   �wh���# S�u�v���YY�E�����   �u��vh����u�Fh=0�tP苮��Y�^hS�=����Fp��   �P���   j�  Y�e� �C����C����C���3��E��}f�LCf�E��@��3��E�=  }�L��P�@��3��E�=   }��  ��X�@���5X�����u�X�=0�tP�ҭ��Y�X�S���E������   �0j�  Y��%���u ��0�tS蜭��Y������    ��e� �E��U���Ã=�� uj��V���Y���   3�Ë�U��SV�5�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�T�t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�T�t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=X�th���   ;�t^9uZ���   ;�t9uP��������   ��  YY���   ;�t9uP�ګ�����   �9�  YY���   �«�����   跫��YY���   ;�tD9u@���   -�   P薫�����   ��   +�P胫�����   +�P�u������   �j��������   =X�t9��   uP蒣  ���   �A���YY�~P�E   ��T�t�;�t9uP����Y9_�t�G;�t9uP����Y���Mu�V�����Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu����tV�s���Y��^�3�_]�jhx��%���������P��Fpt"�~l t�����pl��uj �����Y���8����j�  Y�e� �5����lV�Y���YY�E��E������   �j�  Y�u�Ë�U��E���]Ë�U���(  ��3ŉE�S�]W���tS�{  Y������ jL������j P�|�����������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M���������������j �����������P�����u��u���tS�z  Y�M�_3�[�[����Ë�U��V�5������u����������^]��5�����Ë�Vj� �Vj������V���P���^Ë�U���u�u�u�u�u�����̋�U���5�������t]���u�u�u�u�u�����3�PPPPP��������3�VPPPPP����j� �Vj������ V���P���̋�U��]������U����u�M��v����E����   ~�E�Ph  �u��  ������   �M�H%  �}� t�M��ap��Ë�U��=�� u�E����A%  ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u���  ������   �M�H���}� t�M��ap��Ë�U��=�� u�E����A��]�j �u����YY]Ë�U����u�M��q����E����   ~�E�Pj�u�}�  ������   �M�H���}� t�M��ap��Ë�U��=�� u�E����A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u���  ������   �M�H���}� t�M��ap��Ë�U��=�� u�E����A��]�j �u����YY]Ë�U����u�M��s����E����   ~�E�Ph�   �u�|�  ������   �M�H%�   �}� t�M��ap��Ë�U��=�� u�E����A%�   ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u���  ������   �M�H���}� t�M��ap��Ë�U��=�� u�E����A��]�j �u����YY]Ë�U����u�M��n����E����   ~�E�Pj�u�z�  ������   �M�H���}� t�M��ap��Ë�U��=�� u�E����A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Ph  �u���  ������   �M�H%  �}� t�M��ap��Ë�U��=�� u�E����A%  ]�j �u�~���YY]Ë�U����u�M��i����E����   ~�E�PhW  �u�r�  ������   �M�H%W  �}� t�M��ap��Ë�U��=�� u�E����A%W  ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Ph  �u��  ������   �M�H%  �}� t�M��ap��Ë�U��=�� u�E����A%  ]�j �u�~���YY]Ë�U����u�M��]����E����   ~�E�Pj �u�i�  ������   �M�H�� �}� t�M��ap��Ë�U��=�� u�E����A�� ]�j �u����YY]Ë�U��}�   ���]Ë�U��E��]Ë�U���u�u�9���YY��u�}_t]�3�@]Ë�U���u�o���Y��u�}_t]�3�@]Ë�U���u�u�~���YY��u�}_t]�3�@]Ë�U���EP����Y��u�}_t]�3�@]Ë�U��E�� ]Ë�U���SV�u�M��*����]�   ;�sT�M胹�   ~�E�PjS�,�  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P��  YY��t�Ej�E��]��E� Y��U���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P貏  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=�� u�E�H���w�� ]�j �u�����YY]Ë�U���(��3ŉE�SV�uW�u�}�M��إ���E�P3�SSSSW�E�P�E�P�9�  �E�E�VP�ξ  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�?����Ë�U��j �u�u�F�����]Ë�U���(��3ŉE�SV�uW�u�}�M������E�P3�SSSjW�E�P�E�P�y�  �E�E�VP��  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����Ë�U��j �u�u�E�����]Ë�U���(��3ŉE�SV�uW�u�}�M��Y����E�P3�SSSSW�E�P�E�P��  �E�E�VP��  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������Ë�U��j �u�u�F�����]���������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u�f�����   u������r)��$����Ǻ   ��r����$���$� ���$�����@�d�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I �ԅ̅ą���������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$����� ���(��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�<��I �Ǻ   ��r��+��$����$������Ć��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I @�H�P�X�`�h�p����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�����������ȇ�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��EV�5�������t�i����    ����������^]á��Ë�U��UVW��t�}��u�2���j^�0�������3�E��u����+���@��tOu��u� �����j"Y�����3�_^]Ë�U��MS�YV�u3�;�u�����j^�0�)������   9Ev�U�;�~��@9Ew����j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W�>���@PWV�������3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0��3ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f���  �u܉C�E��E��C�E�P�uV�������$��u�M�_�s^��3�[�"�����3�PPPPP����������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j����YË�U��E�M%����#�V�u������t$��tj j ��  YY�����j^�0�
������P�u��t	�k�  ���b�  YY3�^]Ë�VW3�����<���u�����8h�  �0���0���tF��$|�3�@_^Ã$��� 3����S�<�V���W�>��t�~tW��W�̕���& Y����м|ܾ��_���t	�~uP�Ӄ���м|�^[Ë�U��E�4Ű��|�]��t$j ���h�   �ȸ��Y�jh�������3�G�}�3�9��u����j�3���h�   蔸��YY�u�4���9t���mj����Y��;�u�_����    3��Pj
�X   Y�]�9u+h�  W�0���uW����Y�*����    �]���>�W�Ȕ��Y�E������	   �E������j
����YË�U��EV�4Ű��> uP�#���Y��uj�����Y�6���^]Ë��  Ë�U��E��E�A3��A�A�A]� ��V��~ t��F� �v�F�VY�F�F��u�^Ë`����u3�À�0|��9��/A�`��3�� ��t݀�A|*��P%���A�D¿�`����@uۊA�`���@t���Ë`�SV� @  W3��9_u	A��`��<A|<Z��   <$�1  2�A�`����B��  ��  ����  ��$�T  �yPuAA�`����J�n  �� �[  ��FtHH���L|y��M~��O�I  ��QufA�`��\������A� �  A�`��t��    �����������  ������   ��t
��������#�ȃ�tE��t#��t
���  �  ��t��?����<�������4��t�濁΀   �%��������   ���t�������@������������ �P  HHt*HHtHHu���������   �3  ��������   �"  ��t��������   �  #��  ��/�O�����5��   ��A�=����������� �  �y  ���  ��  A�`��<0|<9���Dѣ`������   �  ���  �9  ���  I�.  �� �  �#  ��C�  H��   H��   �������A�`���<0��   <5��   �� �  ��0�   ��t
����������������t��������   ���������   �t��    ����������� t=HHtHH�1�����t��?����r�������j��t�濁΀   �[��������   �M��t�������@�>��������43Ʉ�������  �  �������� �  ��������� �  ��� |  A�`��U  �<0�,  <8�$  ��A��Ё�����`����y����$���� �  ��t��������   ���������t�������@��   ��������   ��   � �  ��t��������   ���������t�濁΀   �   ��������   �   � �  ��t��������   ���������t��?����w�������o��������e�������� `  �W��������    �I�������� h  �;�������� p  �-�������� x  �<9uA�`����  �3Ʉ�������  ��_^[Å�Œ�6�N�@�\�j�x��p��Ѓ�áp����Ѓ�áp����Ѓ�áp����Ѓ�áp����Ѓ�áp����Ѓ�áp���`3�<`����áp����Ѓ�áp����Ѓ�áp���	�Ѓ�áp�%   áp�%    áp�% @  áp����Ѓ�áp�%   áp����Ѓ�Ë�U��p��Ш�E��hmu��]Ë�U��VW�}������} ��tW�Y�d��uj_�FS;�sE�   ;�w8jh  �@�������t�  �3���t�N��t���F+߉F�^�	3��+ǉF�F�N�D[_^]� ���  �@ �`� ��Ë�U����M���I�H]� 3��y���3�9����AË��H   ËA�����3�9t
�A   t@Ã9 t�I   �3�9t
�A   t@ÁI   ËA����ËA����ÁI   ËA����ÁI    ËA����ÁI @  ËA����ÁI �  Ë	��u3�Ë� �	��u2�Ë�`��U��	��u�E]� �]�`��U����xt�M�Q��~�P]� ��U����M���I�H]� 3��9	��Ë���Ë�� �nË�U����M� �n�H]� 3�@ÊAË�U��E;Es�I�@]� ��U����M� o��t�Q��t��u3ɉH]� �A��t� ��t����"3�ËA��t� ��t����b2�Ë�U��A��t� ��t���]�b�E]� ��U��U���PJ��҃����� o�P]� �AÃy����$ Ë�U��3�A���u]	���o3ң|����������������   ������   ���������   ����E��w
k�|�]ø��]Ë�U����M�H��H�M� o�H]� ��V��~ }�N�SW�~��؋����_�^[�F^Ë�V��N��P��u	�N�^�`^Ë�U��V�u��N�u��P;Es�u�N�P�R^]� 3�8t@A�9 u�Ë�V���t+Ȋ�@Nu�^Ë�U��} u3�]Ê��t:uAB�Mu���
+�]Ë�U��U�����H,�	��d��`��U��tV�u�5l��h�^��%h� �%l� �X��M�p��M�T��t��x� ]� ��U���3ɸ  ��!E�!E�Q�E�Ph�l�E�P�u�M��M��N>  �E���Ë�U����e� �e� �  ��!E�!E�j�E�Ph�l�E�P�u�>  �E���Ë�U���u�@��u�����]Ë�U��EV�uW�}+�;�~����t�E��+ǋ�S��AJu�[�7_^]Ë�U��} V��t0j j�@�������t�u�������3��������$�F��& �F �f� ����^]� ��U��V��M�f� ����t	��t3�����& �F��uQ�����Y���u�F��^]� ��U��S�ًV�uW��t<��u���xVW�@����������t&��}���u�����T>�RV�P�  ���t� _��^[]� ��U��VW�}���t.j j�@�������t��H�� o�H�x�3����u�F_^]� ��U��V��& �F �f� ���} t&j j�@��5�����t�u���D����3����u�F��^]� ��U��EV��f� ���F��uP����Y���u	�F��& ��^]� ��U��V��>	t6W�}�? t,j j�@�������t���O�H�3���t���D�_��^]� ��U��E��	w1����t;��L���E��I�H� �E�`� ���  �@��Mj������E]� ��U��VW�}���(o��t1�} t+j W�@������F�~��t��t�M+Ȋ�@Ou���f �f _��^]� �AËA��t�I�D��2�Ë�U���q�q�u�u�������]� ��U��yujh4o�u�u���������E]� ��U��`��8@�uu�M�`�������
�u�bI  YY�E]Ë�U���u������EY]Ë�U��V��~-�> �Et��t��t��tP�����YP���q����P�������^]� ��U��SV��3�9t�f� ���F��_W�};�tR�E;�tK+�tAHS�@�tj�����;�t%�u��W�w����j����;�t�� �n�H�3��;�u
�F��F_^[]� ��U��3�V��F�f� ���8Etj�EP�W�����^]� ��U��E3�V��V�f� ���;�t3�8tA8u�;�v	QP��������^]� ��U��V�u3�W���W�g� ����;���   8��   �E��:EtK<_t<<$t8<<t4<>t0<-t,<a|<z~$<A|<Z~<0|<9~<�r<�v�p�   t;BA����8 u�R�u����������t@�:Mt�' �G�� u
�G��G��_^]� ��U���$��3ŉE�S3�V��W�F�f� ���}���E�j j
�uO�u�`�  ��0�E]���UuލE�+�PW��������M�_��^3�[�J~���� ��U���(��3ŉE��EV��3ɈN�f� ��W�}���M��M�;�|9Ms�U����E��؉US�3�Qj
P�uO���  ��0�E��M��ȉ]�u�[8M�tO�-�E�+�PW���]����M�_��3�^�}���� ��U��V�u�u��A�ΉF�������^]� ��U��V��~.�E���u�@P���������> u
��@�F�Q���M�����^]� ��U��W���RV�u��tI�? uV�m����<�F��t<t��P�k����&j j�@�������t
V�������3�P�������^��_]� ��U��3�V��F�f� ���8Etj�EP�W�����^]� ��U��E3�V��V�f� ���3�8tA8u�QP���"�����^]� ��U��QQ�`�� ����   ����A�`���w�U��e� �� ��jYщU��p�������tK����� t0+�t)+�t!+�t+�t��t+�u*j�j�j�j�	j�Q�j�{�����P�M��5����E�M���M��H�ËE�`� ���  �@�ËMj�����E�Ë�U��`�� ��t,<At�E�`� ���  �@]ËM�`�h<o������
�Mj������E]Ë�U��V�u�u��A�ΉF�������^]� ��U��V�u�u��A�ΉF�������^]� ��U��V��~=S�]��t4�> uS�"����'j j�@�������t� �n�X�3�P�������[��^]� ��U��W���OSV�u3�;�tB8t>9uV������2Sj�@��A���;�t3�8tB82u�RV��������3�P���u���^[��_]� ��U���S3�V�u�^�f� ���E�   �8^��   W�`�� <@��   <Z��   9]�t�]��	j,��������=`��:���   ����0��	w!�T�P�E�GP�=`������P���S����Y�e�  ���E�P�E�P�]��@  �`�+�YY��~�T��9	t	�E�P�m����E�P������9=`�u�f� ���F�8^�8����	j�������_��^[�Ë�U��QQ�E�V�u��@hDo�ΉF�r����E�P�j,  YP������j}�������`��8@u�`���^�Ë�U��QQ�u�M��u�u�����������E�Ë�U��QQ�u�M��u�u�2������e����E�Ë�U��QQ�u�M��u�u� ������A����E�Ë�U��V�u�u��A�ΉF�g�����^]� ��U��V�u�u��A�ΉF������^]� ��U��`���S3ۀ9QuA�Lo�`����u�Mj�����E�	  <0|L<9H���/�AR�`�P��t�M��J���P�E�SP�+�������M��2�����M��@�A���   VW3�3��)��tI<A|2<P.������A�����A���`��<@uӊA�`�<@t"�E�`� ���  �@�b�Mj������E�S�} WVt��t
�M�������M��
����$��t�M�����P�E�SP�o�������M��v�����M��@�A��_^[�Ë�U����`�� �e� �e�  ������   ����Ѓ�w|�$�ϧh�o�h�o�h�o�hxo�M������`�� �`���1tHHtHHtHHu$�E�P�E�Phlo�M�������������M��U���U��M��E��P�ËE�`� ���  �@�ËMj�����E�Ð7�7�>�>�Y�E�L�L���U��`�� ����X��   HH��   �E�P����Y�M���uh�`�� ��t]<@tS<Zt�E�`� ���  �@�áp��`����Ш��ou��oP�E�P�M��'�����M��@�A�����`��E�U���H�áp��`����Ш��ou��oP��`�h�o�M�����E�Ë�U��`�� ����tL<Zu�`��U��E3Ɂ�  ����P�ÍE�P�����YP�E�Ph�o�M��L���������j)�u�M��!j)�u�E�jPh�o�M��#������!������!����E�Ë�U���$�e�  ��S3�3��`��`����V����AW�� ���a  N�*  N�  :��  �`��R:���   9]t�E�`� ���@�L  �`��������t�Ѓ�vA�e� ����e�� ��j�E�P�M��E�,�]�����SV�M��R���P�E�P�M�������@��E��M�j>�M�E������`��:$�E�M��E�M�u�`���M�j^�M�E������E�E�E��E��`�8t�`��
j�M�������M��E�U�� @  ��H�v�Mj������E�g�E� �l�K9]������E�e� ���!}�� j�E�P�M��E�>�]�������9]u�M��8&��lt�pl��E�`��X!x�_^[�Ë�U��`���8S3�8�B  �K����E�;�}�]�9]�u�E�j]P�E��M��  �e�  ��VW�}�   �]��wtfh�l�M�������W�E��M���tS�`�8tJ�E�SP����YYP�E�Pj[�M�������������E��E�E�j]�M�E��(����E�P�M������}�~�9tn�wt�E�P�E�P��������M��@�MW�E�Pj(�M��(����������E��E��E�j)�M��E�������E��E�E��E�E�P�M��I����E�E��E�E�E�P�E�P�8  �E�U�YY�M��_��H^�   �E9t`P�E�Pj(�M������������E؉E�E�h�o�M�E������E�E��E�j�M��E������E��E��E�j]�M��E������E��$�E�j]P�EЍM�jPj[�D������o������o���P�u�<4  �EYY[�Ë�U����E�j P����YYP�E�Pj`�M��������o���j'�u�M��&����E�Ë�U��j�u�Z����EYY]Ë�U��j �u�D����EYY]Ë�U��j �u�.����EYY]Ë�U��E��� SV�u3ۉ�@C�F:��4  �`��9 �  �E�P�����E�Y�E��E�j �M��E�����V�E�P�M��������@�F:���   �`��8@��   hDo�o�`�� ��tp<@tl�E�P�#  YP�E�Pj`�M���������d����E��E��E�j'�M��E������E�P���$����`��8@u@�`�8^6�8@th�o������8^~�8^�`��8 uS�������j}���@����`��8@u,�`��$:� V�E�PS�M�������������E���E�F��^[�Ë�U����u�M��a����`�� �`�<@u|�`�� �`�<_uk�`��E�j P�����E�j P�w����`������t��@t@�`����u�8 u�MHj�`�������E�ËM�@�`��E��M��H�ËE�`� ���  �@�Ë�U��QQ�`�� ��u�Mj�����/j <?u�`��E�P�����Pj-�u�#������
�u�����YY�E�Ë�U����   ��3ŉE��`�S��`�V�uW����D�#  �u  �� �   ��0��   O��   Ou@�E�P�O�����x���P�C����}�YY��   ��|�����   jd�E�P�M��0�����u�f� ���& �F�6  �E��E�<-u�E��E��E�.��E�.��x���PVje��`���P�E�P��@����������������������  �`��8@u�`�h�o���]�����  ��8���P��  YPVh�l��p����9����V�p����  �`�j���+����  ��E�x  �0�����J��   ��Qt;��R����j ��x���j P�  �E�P������x������|������F�0  �E�P������p� @  Yt*j�E�P�M�������E�P��  P�t�YY��tP�����E�P��x����M�P��Du'h�o�c���������h�oV��x����{����   hLo��j{�M�������H|%��J ��P���P�  YP�M��>���j,�M�������Ft,Ot	OtFOt#OuV��h���P�-���YP�M�����j,�M��j�����X���P����YP�M������j,�M��J�����H���P�����YP�M������j}V�M������V�  Y�M�_��^3�[�1k���Ë�U��`�3Ƀ�8��   9Mt7�8Xu2@�`��E9u�Mh�o�D����   Php�u�����   �8Yu�u@�u�`������YY�uV�u�E�VP��-  �FYY^� @  t$�E�P�E�Php�M���������#����U��M���    t�E�P�E�Ph�o�ӋM��U��E��H���uj�u�d������E�Ë�U���u�u�����EYY]Ë�U���|��3ŉE�S3�V�u�^�f� ����y��E�   8^��  W�  ���`��:���  ��@��  9]�t�]��j,�������`���ʃ�0��	w@�`�Q�\��E�P�����M  !}�E��]��Xu@�`�h�o�M�������  ��$u@8t�`��E�P�:�����   ��?��   �E�P������p� @  Ytgj�E�P�M�������E�P蚿  P�t�YY;�tP됍E�P�E�Ph�o�M��I����������E��E؋E�h�o�M؉E������E؉E�E��]�E�P�E�Ph�o�M��	������J����E��EЋE�h�o�MЉE�������EЉE�E��!}čE�P�E�P�]��p/  YY��@�M�E�`�+E���~�\��9	t	�E�P�����E�P������8^�J���_�M���^�y�3�[�$h���Ë�U���   �`��S3۹  ��!M�!M�V3�@�]��]�`���A��  �g  ;��]  ��/�J  ��1~[��9�<  �@��4��l�M�����9]�t(�E�P�E�Ph�l�M���������(����E؉E��E܉E��M��E��M��H^[��!M�]�8]t|��x���P�*���YP�E�Pj<�M��n�����������E�P�M������M�;�t��P<>u
j �M������j>�M�������E;�t� �`�8u�M��E��M��x���@�`�S����p���SP��  ��@���M��E��5`�;�t+�~�1u%�E�P�E�Pj~�M���������<����M��E�M��E�9]������E�P�M�����������H�`��Mj������E�������B��  ��  ��Z��  ��_��  �@�`���O��   ��D��  ��9kt@;�t���/��  ��6~��8��  �@��4�`m�M�E�����@��4�`m�*����@��4�`m�M�� ����M�� �  �U��E��A�����?t9��@�$  ��B�  ��C�  jh�k�E�P�f����M����   ��@�`�;��������0��  Shp�ǃ�T��  ��S��  ��P��  I�����I��  �@��4�Dm�M��n����`�� :�uj�u�M��[�����������0�m  ���d  �4��n�M��-����`�� �`���0��   ��1t��΃��B  �`��2����E��E�E��E�E�P�M�����j,�E�P�E�P����Y�������P�M������j,�E�P�E�P�����Y������P�M������j,�E�P�E�P�����Y������P�M�����j)�E�P�E�SP�����YY���u���P�M�����j'�u�M��_��������E�SP�,  �E�YY�E�E�j �M�E������E�E��E�E�E�P�M��=����M��O�@��4�Dm�M������S�E�SP������@���M��E�;�t�   t�E�`� ���@�������M��E�P�u������������U|҃�V��   ��W~ă�Y��   ��_u��@�`���A|���D~
��F~��J��@��4��m�����@��4��m�M��N����`��8?u%�E�P�  YP�M��Z����`��8@u�`���E�P��  YP�M��5���hp�M�������M�E��M��&����@��4�Dm�����@��4�Dm�����3�F�@��4��l�M�����;������9]�������M�   �������U��`���   �8?�+  �x$�!  �M���M����X����S�\�V�5T��M��T��M�W�=X��X�����X����`��\��8?�E� u@�`��E�P�E�jP�����j�E�jP�   ��@���E��M��u�x��}� uf�E�P�Y���YP�E�Pj<�M������������E�P�M�������M��t��P<>u
j �M��-���j>�M��#����} t�`��8 t�`��E�M�=X�_�5T���M�^�\��H[�ËE�`� ���  �@�Ë�U���8��3ŉE�S�`����V�u��0�uȃ�	w�X�PCV�`����������  �e� W�  ��!}��?uJ�E�j P�D���YY��@�E�`��M�@�`���@�W  H3ɣ`�8��AQ�M�������;  �Hp�����E�   ���t:uAF�M�u��	�+�u���`��0�8pj�ˋ�[���t	:uAFKu��	�+���   �`����E�P�o����p� @  Yt2j�E�P�M��h����E�P�8�  P�t�YY�M��tP������   �M�h4p������E�P�E�PV�M�������������EԉE܋E�h�o�M܉E������E�P�M�������?�} t�`��8@u�M�3�#��`��E�M��j@h`��M�������@�M�E�} _t�X��9	t	�E�P������M�Eȉ�M�H�M�^3�[��^���Ë�U���SV�uW3�S�E�j�^�� ��!~P���������@���F:�u?�`�� :�t4<@t;V�E�Ph\p�E�P�E�P�  Y����������������@�F�`�� <@u�`��N:�t!~�F��?9uj��������0V�E�Ph\p�E�Pj�M��{������������������@�F_��^[�Ë�U���u�����EY]Ë�U��p��� VW����3���G#�t�   t3��`�� �e� �  ��!u��`��� ��   ��Tt^HtTHtJHtHt
Hu\h�p�Mh�p�F�E�P���_���YP�E�Ph�p�M�������������E��E��E�E��h�p�hxp�hpp�M������e� !u��t�E��E��E��E�E�P�3���Y�E�P�M��~����M��E��M�H��M�`�hap�2����E_^�Ë�U��`��8?u'@�8$uj�u�p���YY�"j j �u�`������j j�u�������E]Ë�U���j ������P�M�������`��8 tP�@�`�����0t1HHt��uA�E�`� ���  �@�ÍE�P�X���YP�M������h�o�M��P����
j�M��p���h�p�M��7����M��E��M��H�Ë�U���XSVW3��  ��!u�}������M��99t�A   �E�   u�}����  u�E�`� ���@�8�_  ����  uQj�u�������E�A  ����  u��E��I�'  �]��e� �  �   �   �M  3��]�!}�}�   ���E�����t%   �#���t��%   ;��  �}� ��t%   �#���t��%   =   ��  =   ��  �� @  t_�p���������t7���Шt.�E�P�,���YP�E�Pj �M���������>����E��E��E��E���E�P�����YP�M�������   �U��Å�t%   �#����,  9}��#  �E�j P�����YY�M�E�P�E�Pj{�E�P�����������P�M������E�P�n����   Y�5p�u>�E�P�E�Pj,�M��$����������E��E��E�h�q�M��E������E�P�M��N���h�q�M�������E�P�D����p�Y���������/  ���������  ���  �E�P�E�Pj �M������������E��E��E�j �M��E��C����E��E��E��EčE�P�M�������M��EĉM��E���  !u�!u�!u�!u�!u�3��}��}��}��}؉}Ћ�;�t%   �#�;���   ;�tw��%   =   u>�E�jP�����EȉE��ẺEčE�jP�s����EȉE��ẺE��E�jP�\������;�t'��%   =   u�E�jP�:���YY�EȉE��ẺE�E�jP�!����EȉE؋E�YY�E�3�9}�tF�}� t��%   =   t2�p���`<`�E�Pt�����Y��@�MЉE������YP�M��c����p���������t/���Шt&�E�P�E�P�E�P�}���Y��������M��@�E���E�P�_���YP�M������E�8 tA�}� t0�p�   u$P�E�Pj �M���������8����E�P�M��������@�M��E�!u�3��}�9}�tE�E�WP����YYP�E�Ph�q�M�������������E�P�M�������p�   tA�M���  3�Wj�@������;�t�8�@ �`� �����E�WP�#���YY��@�MȉE̋u��Å�t%   �%   ���  ����   ��%   =   uz�E�P�E�Ph�q�M��������E����E�E��E�j,�M��E��w����E��E�EĉE�E�P�M�������E�E��E�j,�M��E��I����E��E��E��EčE�P�M�������.��tN��%   =   u@�E�P�E�Ph�q�M��x����������E��E��E�j,�M��E�������E�P�M��x����h�q�M��"����E؉E��E�h�q�M��E��	����E�P�M��D����E�P����YP�E�Pj(�M���������C����E��E��E�j)�M��E��u����E�P�M�������t��%   =   t�E�P�M�������p����Ш�E�Pt�
���YP�M������������YP�M��z����p����Ш��  ����  �E��Mȉ�E�G�ẺM��E��  �u�M��q����E�� |  ����   ��#с� h  u�E�P�u�M���YY�@�������   ��#с� p  tم�u|��#с� `  uOP�E�P�?����E�YY�E��E�j{�M��E��c����E��E��E��EčE�P�M������h�q�u�M�������������u��#�;�u�E�P�u������i�����t��#�-   ���% `  ���@���   ��t%   �#ƅ�t$�E��Ӂ�   +����B�����t
hdq�   �}� ��t	#�-   �% `  ���@����t%   �#ƅ�t%�E��Ӂ�   ��   ���B�����th0q�Q�}� ��t	#�-   �% `  ���@����t%   �#ƅ�t-�E��Ӂ�   ��   ���B�����th q�M��h�����}� u��#�= x  ������}� t��#�-   ���% `  ���@����t%   �#ƅ�tX�M���%   3�=   ����Ʌ�u�M�3�=   ����Ʌ�t'�E�P�E�Ph�q�M���������:����M��E��R����E�P�E�P��  YY��M��@�9����M�   3Ҿ   ��9U�t#�+��% `  ���@;��s  �p���	�Ш�M  ��9U�t#�+��% `  ���@;�tG9U�t��%   -   ���@�3�@;�t(�E�P�E�Ph�p�M��<������}����M��E��M��E�U���t��%   =   ��   ��t��#�+����% `  ���@����t%   �%   ����   �Å�t#�+��% `  ���@��t��%   =   tP�Å�t#�+��% `  ���@��t��%   =   t(�Å�t#�+��% `  ���@��t6��%   =   u(�E�P�E�Ph�p�M��Q����������M��E��M��E�p����Ш�  �}� ��t#�+��% `  ���@��t4�}� ��t$�3�<@���	#�+����@��t�E�P�E�Ph�p�   �}� ��t#�+��% `  ���@��t4�}� ��t$�3�<����#�-   ���@��t�E�P�E�Ph�p�G�}� ��t#�+��% `  ���@��tF�}� tj ���X���	��#����@��t(�E�P�E�Ph�p�M��=������~����M��E��M��E�}� ��t#�+��% `  ���@����t%   �%   ��t4�p�   u(�E�P�E�Ph�p�M�������������M��E��M��E���   t%�E�P�E�Ph�p�M�������������E��M��E�E��M�H_^[�Ë�U���$SV�    W�5p�t0�%p������E�j P�  	5p�YY�M܋E��M��H�!  �`����?�   @�`�8u#8Hu�E�P�����`�Y�@�`��8 u�밍E�P������u�]�3�@Y��t��   t�E���e� ����#�:�~�E�0�X�  �`�� ����   <@��   �E�P�  �E�Y����   �=x� ��   �E�P�M��x� �u�]������`��8@�u�]�u�]���   �E�P�4  ��M�H�M���@�M�M�E��$\p�����E�E܋E�E��E�P�M��=����u܋]��4�E܋E�h\p�M܉E�������E܉E�E��E�E�P�M������u�]�]��u�}� t��t	��   �]�� �  ��tډ]���������   ��������`�� ��t<@t�E�`� ���  �@�X�`��p�t)�}� u#��u�e� �e�  ���E�P�E�P����YY�p����E�P�u�����YY���u��Mj�3����E_^[�Ë�U���   SV�u3�W�� ���^!~��]�&  �`�� :��   <@�  8x�t8y��]  9tSV�E�Ph\p��p���������������E���E�F8]t'V�E�Pj[��h����[�����������E؉�E܉F�]�`��9?�p  A�`����$�I  H��   ��t^HH��   ��Vt��X���P��H���P�����Y�>  �E�Pj]�E�PS�E�AjP�`����������������8����E�  �A�8_uK�y?uE�`�V��P���PS�E�SP�O���������������@�F�`��8@��   �`���   ��`���P�����YP�E�Pj`�M��K����������E�E��E�j'�M��E������V�E�P�M��sj@h`��M�����V�E�Php�M��0������q����E���E�F�X��9	tD�E�P�����9��x���VIP�`��E���E�VP�E�SjP���������!������@�F8^������`�� :�t<@tJ!~�F��?9uj��������0V�E�Ph\p�E�Pj�M��������������������@�F_��^[�Ë�U��`����8��u�uj�u�
����E���À�6|��9~��_t�E�`� ���  �@��S�ك�6@�`���)u4���t�ك�=@�`���|&����uj�u�����E���L  ��x��~������u�E�`� ���  �@�%  �e� �e�  ��V�u�W�E��F�����E���   �E�P�E�Ph\p�M��t����������E�E��E�E��`��8 tC�E�P�1���YP�E�Pj �M������������E��E�E�E�E�P�M��H����E�E��E��"�E�P�E�Pj�M��������C����E��E��E�E��`�� ����   <@��   �p��`���`<`�E�Ptq�����Y��@�M��E�����   �p����Ш�E�P��   ����YP�E�Pj �M��Q����������E��E�E�E�E�P�M������E�E��E�E��S����YP�M��3���돋E�`� ���  �@�  �E�P�u�M�j�'������Z����~  �'���YP�M������p����Шt&�E�P�E�P�E�P����Y��� �����@�M��E���E�P�����YP�M�詿��3�9t;�E�P�E�Pj(�M��s�����������E��E�E�j)�M�E������E�E��E�E�Sj�@��ý��;�t�X�`� ������3��E�VP�����E�P�������P�E�Pj(�M��������p����E��E�E�j)�M�E������E�P�M��/����p���`<`t;�t�E�P�M������p����Ш�E�Pt�9���YP�M��������(���YP�M�詾��;�t�E���E��F�M؋E��M܉H��Mj�����E_^[�Ë�U���T�`�� SV�  ��!u�W3��E� ����  <$u.�u�E�P�EP�E�P�7����Mԃ�;�t�E��M؉H�@  �`��3�<A��!u��؉}�J��+��+�3�!u�U�Ã���   HtN���n  �p����Ш��   ��t)�E�j �MԉUԉE��U���j	�������P�E��M��   j	�   �p����Ш��   ��t7�E�j �M܉}܉E�����j
賻����P�E�P�M������8�@�}�E��j
菻����P�M��I����}��g�p���������tW���ШtN��t7�E�j �M�U�E�����j�G�����P�E��M�P�-�����@�M�E��j�#�����P�M�������`��`��8$u�u�E�P�EP�E�P�����M̃���u#�`��3�<A����J��+��+ڋU������E��M��J����9 tA�`�����   �uV�M��^���3��E܋EȉE��E�P�M��p����}� �E܋M��E�M�t4�M�j �M܉E������E܉EԋE��E؍E�P�M��6����EԉE�E؉E���t7�E�j �Mԉ}ԉE��z����EԉE܋E؉E��E�P�M�������E܉E�E��E�����   �} t�E�`� ���  �@�  �> tx�E�P�E�Ph\p�M�������������EĉE�EȉE��`��8 �E�Pt�E�P�E�P�<���Y��������@�M���E�Pj�M��G������z����EĉE�EȉE���`��8 t�E�P�����YP�M�������`�� ��uj�M�� �����`�<@�+����p����Ш��t7��<uJ�} �����E�P�E�P�E�P�����Y���������@�M�E����<u�E�P����YP�M��s�����t(�E�P�E�Ph�q�M��h����������EĉE�EȉE���t(�E�P�E�Ph�q�M��;������|����EĉE�EȉE�3һ   9U��   �u9t`�N��uB�E9t;P�E�Pj �M���������5����EĉEԋE�j �MԉE��g���V�E�P�M������7��   t��E���E��,V��E9t"P�E�Pj �M��n�����������E�P�M������M�ˀ}� t��    �E�U��5���9}uk�u9>tZ�F   uA�E98t:P�E�Pj�M��M����������EĉEԋE�j �MԉE�����V�u�M��^����$Vj�u���������E98tP��Mj������E_^[�Ë�U��� �E��  ��!U�3�!M�#d���tq�:?u]�B<@u2�`��E�P����YP�E�Ph�q�M�������������M��E��3<$u �E�j P�����YY��@<u�d��`��E�P�����Y��@<u3���<t�p�   u�`��: u�M��E���5d��M������h���u(�M���t��@�l������P�@�Y�h���t>�5l��M�P�-����h������ u@�
B�@�8 t���
B@���u����h��Ë�U��QQ�`�� S3�V:���   <6|<9~<_uN�u�M��x����E�u9t9t	�F   u	P�M�����9t	V�M��t����E�P�u�����YY�E�   �uS�u�E�V�uP����3��>*��P�E�P�u������ ��j�M������u�M�������u9t	V�M�����W�}9t9t
j �M��\���W�M�������M��E��M��H_^[�Ë�U��h�l�u�u�u������E��]Ë�U��h�l�u�u�u������E��]Ë�U���u�u�u�u�����E��]�jdh���p���}3�;�u3��rj����Y��t�j�ƭ��Y�u��=@��E�D��5P��5H��5L��EPV�u�u�u�M��v����M�������E�@��έ���E������	   �E���o���j�i���Y�jdhا�o���}3�;�u3��rj�v���Y��t�j�,���Y�u��=@��E�D��5P��5H��5L��u �u�u�u�u�M��ܷ���M��a����E�@��4����E������	   �E��Do���j�ϫ��YË�U��`�� ��$SVW���l  �`��e� ���  ��!u��ǃ���E� ��NR�-  ��C��
�  ����$���h|r��  htr��  hpr��  hhr��  h`r�  ��O��  ��  ��S��  ��X��  ��_��  �`�� �`��E�����M��   ��L��   ��Ge��F}V��t=��$t�������   hXr�C  �u�E�P�����PhPr�u��������m  �`�j�M��,����H  hHr�  ��H|x��I~��Knh@r��   h8r��   h,r��   ��N��   ��OtW��RtK��Wt?�����w0�E��`�P�?����PY��M�U�����   �E��P��  h$r�~hr�whr�pj�[�E��e� !u��M�H�M�����4  h�l�E�P�E�P�E�   	u�P�\������u�uh�l�M��ҿ���M�E��M���   hr�h�o�M��̽���2�߃��"�E��5���hxo�M�讽��h r�M�胿������W����ǃ�Ct@jY+�t*+�t&+�t"+�t��uP�E���Et+�t+�t+�t+�u7�E�P�E�Phlo��E�P�E�Ph�q�M��<������}����E�E�E�E��E�8 t"P�E�Pj �M��������S����E�P�M��(����M�E��M��H�j�8 u8��t!h�q�M��ؼ����t!h�q�M�訾�����th�q�M�貼��h�l�E�P�E�P�u���������uj�u�O������E_^[�Ë�������������   ��U����`�� S3۹  ��!M�+�V�]��s  ��$tj���ut.HtV�u�����YY�c  h�q�M�����9t
j �M�艽��h�l��v�`��E��E�P�E�P�u��   �u��$������  �`��@<$t:���   �E�`� ���@���   �`��`�� �u��Qp��   +�tc��AtJHt4Hu��`�!M�S�E�Ph�l�E�VP�]������P�u�)������   �`�jV�u�����x�`�V�u���������V�W��Rt*HtH�U����M�`�h�r�����@�`��5���h�q�M��ٺ��9t
j �M��[���hhl������uj�u�x������E^[�Ë�U����u�M��R����`�� 3�:���   <?tG<Xt�E�P�u����YY�   �`�9M�u�Mh�o�S����q�E�P�u�M�hp�=����T�`��e�  ��Q�E�Ph�l�E�P�E�P�M�������M��@�E��E�P�u��������E�P�u�M�j��������(����E�Ë�U���Vj j�@�������t�  �@ �`� �����3�V�u������E�P蔱���E����E��E�j �M��E������u�E�P�M�躺�����@�F�E^�����������SVW�T$�D$�L$URPQQh��d�5    ��3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C��&  �   �C��&  �d�    ��_^[ËL$�A   �   t3�D$�H3��Y5��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�?&  3�3�3�3�3���U��SVWj RhF�Q�V _^[]�U�l$RQ�t$������]� ��U��E������������]�jh���f��3�W�u���Y�}�9}u����5������E��E�   �����5������E��E�   ;�t��t�hU����E������   9}�u3��3�W����YÃ}�t�u��U�Y3�@�lf��� ��U��E��cV9Pt��k�u��;�r�k�M^;�s9Pt3�]��5��������V����d���V����`�jh���e���e� �u�]����  ����  j_;���   ����   ����   ����   ����   ��t��t	����  ��U��������  �@c9~\u'�5�c�Y��Y�F\���t  �5�cWP�-�����v\�������Y���Q  �H�M�M���.  ����H����ck�V\�x�;��  9t��  j 薢��Y�e� ;�t��u>�=�� u5jh�����3�A;�u�����gi���������E�   �u��+�ty��t��	tN��t(H��   �5������E�;�toV�������a�5������E�;�tNV�������@�5������E�;�t-V��������5������E�;�tV�������E������   �}� u�E��8�]j 蚠��YÃ�t$��t��t��~��~�ah���    跍�������c���j h8��c��3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC��S�����}؅�u����T  �������U�w\������Y�p��Q�Ã�t2��t!Ht��g���    �(���빾�������������
�������E�   P����E�3��}���   9E�uj�s[��9E�tP�y���Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,��c�M܋�c�c9M�}�M�k��W\�D�E����UQ����E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��1b��Ë�U���$��3ŉE��ES�E��EVW�E���P���e� �=�� �E�u}h�r����؅��  �= �h�rS�ׅ���   �5��P��h�rS�����P��h�rS�����P��h�rS�����P�֣����th�rS��P�֣������M�5��;�tG9��t?P���5�����֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3���;E�t)P�օ�t"�ЉE��t���;E�tP�օ�t�u��ЉE��5���օ�t�u�u��u��u����3��M�_^3�[�Z.���Ë�U��V�uW��t�}��u�$e��j^�0�{�����_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f���d��j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�d��j^�0�������݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f��d��j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u��c��j^�0������_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f��c��j"Y���뼋�U��M��x��~��u���]á�����]��Oc���    襈�����]Ë�U��E� �]Ë�U��ES3�VW9]u;�u9]u3�_^[]�;�t�};�w��b��j^�0�U�������9]u��ҋU;�u��ك}���u��+�
�B:�t"Ou����+���A:�tOt�Mu�9]u�;�u��}�u�MjP�\�X�x�����b��j"Y���낋�U��E��t�M���]Ë�U��E��t���8��  uP��/��Y]Ë�U�����3ŉE��E� �@SVW�=��3�VV�u�E��u�׋ȉM�;�u3��   ~Ej�3�X���r9�D	=   w���  ��;�t����  ���P��.��Y;�t	� ��  �����3�;�t��u�S�u�u�ׅ�t VV9uuVV��u�uj�SV�u��H���S����Y�ƍe�_^[�M�3��*���Ë�U����u�M��4���u�E��u�u�uP��������}� t�M��ap��Ã%X� Ë�U��M��tj�3�X��;Es�a���    3�]��MV���uF3����wVj�5�������u2�=�� tV��a��Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u�-��Y]�V�u��u�u�4.��Y3��MW�0��uFV�uj �5���������u^9��t@V�a��Y��t���v�V�oa��Y�8`���    3�_^]��'`�������P��_��Y����`�������P�_��Y����ʋ�U��MS3�;�vj�3�X��;Es��_���    3��A�MVW��9]t�u�F_��Y��V�u������YY��t;�s+�Vj �S��"������_^[]Ë�U��E���]Ë�U��QV�5��������E��u�\_��j^�0賄�����   �  W����   h$s����E���u�(_��j^�0�������   hsP� �����u(� _���5������P�^��Y��I�����P�^��Y�LSV������I��Wh�������;�[t	�u����j�u�օ�u�^���    �^��� �3�_^���������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�hX�h�Pd�    P��SVW��1E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����u�M��S0���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �u�u������]Ë�U��jj �uj ������]Ë�U��jj �u�u�h�����]Ë�U��jj �uj �P�����]Ë�U��jj �u�u�7�����]Ë�U��jj �uj ������]Ë�U��jh  �u�u������]Ë�U��jh  �uj �������]Ë�U��jh  �u�u�������]Ë�U��jh  �uj ������]Ë�U��jh  �u�u������]Ë�U��jh  �uj �z�����]Ë�U��jhW  �u�u�^�����]Ë�U��jhW  �uj �C�����]Ë�U��jj�u�u�*�����]Ë�U��jj�uj ������]Ë�U��jj �u�u�������]Ë�U��jj �uj �������]Ë�U��jj �u�u�������]Ë�U��jj �uj ������]Ë�U����u�M���-���E��t*�x�  u!jj �u�u�y������}� t�M��ap��À}� t�E��`p�3��Ë�U��j �u����YY]Ë�U��QV�uV�7�  �E�FY��u�VZ��� 	   �N ����/  �@t�;Z��� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,��  �� ;�t��  ��@;�u�u裃  Y��uV�O�  Y�F  W��   �F�>�H��N+�I�N;�~WP�u�K�  ���E��M�� �F����y�M���t���t���������������@��@ tjSSQ�z  #����t%�F�M��3�GW�EP�u�܁  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U��Q�C@V����E�t�{ u�E�>�' �} ~0�E� �M���n����E�>�u�?*u�˰?�X����} Ճ? u�E��^�Ë�U��E� � �@�]Ë�U��E� ��A��Q�]Ë�U��E� � f�@�]Ë�U���  ��3ŉE�S�]V�u3�W�}�u��������������������������������������������������������������*���W����������u+�W���    ��|�������� t
�������`p�����7  �F@u^V�A�  Y�@����t���t�ȃ��������������A$u����t���t�ȃ������������@$��q���3�;��g��������������������������������
  C3�������9������y
  �B�<Xw����8s���3����Xsj��Y������;�� 
  �$�����������������������������������������������	  �� tJ��t6��t%HHt����	  �������	  �������	  �������	  �������   �	  �������	  ��*u,����������������;��l	  �������������Z	  ������k�
�ʍDЉ������?	  �������4	  ��*u&����������������;��	  ��������		  ������k�
�ʍDЉ�������  ��ItU��htD��lt��w��  ������   ��  �;luC������   �������  �������  ������ �  �<6u�{4u�������� �  �������p  <3u�{2u������������������N  <d�F  <i�>  <o�6  <u�.  <x�&  <X�  ������!�����������P��P� 6  Y��������Yt"�������������V����C��������������������������4����  ��d��  �X  ��S��   tL��AtHHt$HHtHH��  �� ǅ����   �������V  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ��u�Լ������������ǅ����   ��  ��X�"  HHt+���  HH��  ��������������  ������t0�G�Ph   ������P������P�Ł  ����tǅ����   ��G�������ǅ����   �������������|  �����������t;�H��t4������   � ������t�+���ǅ����   �7  !������,  �м������P�v���Y�  ��p�=  �%  ��e�  ��g��   ��it|��nt.��o��  �������������ǅ����   tl������   �`�������������p��T  ���b��������� tf������f���������ǅ����   �>  ������������@ǅ����
   �������� �  ��  ��W���  ������������@�������   ������������9�����}ǅ����   �ju��gucǅ����   �W9�����~�������������   ~=��������]  V��@��������Y��������t���������������
ǅ�����   ��5�����������G�������������P��������������������P������������SP�5 ����Ћ���������   t������ u������PS�5,�����YY������gu��u������PS�5(�����YY�;-u������   C������S�����ǅ����   �������*��s�n���HH�X�������  ������ǅ����'   �������ǅ����   �2���������Qƅ����0������ǅ����   ������   �������� t��������@t�G���G����G���@t��3҉�������@t��|��s����ځ�����   ������ �  ����u3�9�����}ǅ����   ���������   9�����~���������u!������u����������������t-�������RPWS�n  ��0�������؋���9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t����u�+��������(��u�м�������������I�8 t@��u�+����������������� ��  ��������@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����+�������������u%���������������� O������������t���������������������������P�����������������YYt.������u%��������������˰0O�s����������t��ヽ���� ������tu��~q�������������������Pj�E�P������P����{  ����u69�����t.�������������������E�P�������Q��������� YYu��#��������������P�������������#���YY������ |2������t)�������������������� O�����������t��߃����� t�������>�������� Y���������������t���������������r��������� t
�������`p��������M�_^3�[�R���Ðd c�����=�H���� ��S��QQ�����U�k�l$���   ��3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|�����}  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�I}  ��h��  ��x�����  �>YYt�=X� uV�˂  Y��u�6�>  Y�M�_3�^������]��[Ë��` � �s�@ Ë�U����M� �s�	�H�@ ]� �A��u��sË�U��} W��t-V�u�u}���pV���YY�G��t�uVP�~�����G^_]� ��V��~ t	�v����Y�f �F ^Ë�U��EV��f ��s�F �0������^]� ��U��V�uW��;�t�����~ t�v���V�����F�G��_^]� ��s�{�����U��V�EP��������s��^]� ��s�R�����U��V�EP���_�����s��^]� ��s�)�����U��V�u���������s��^]� ��s������U��V����s������EtV�n��Y��^]� ��U��V�u��f ��s�F ������^]� ��U��V����s�����EtV��m��Y��^]� ��U��V�u��������s��^]� ��U��V����s�^����EtV�~m��Y��^]� ��U��V�u���`�����s��^]� ��U��V����s�����EtV�:m��Y��^]� ��U��V�u��������s��^]� Pd�5    �D$+d$SVW�(���3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(���3�P�e��u��E������E�d�    �Pd�5    �D$+d$SVW�(���3�P�E��u��E������E�d�    �Pd�5    �D$+d$SVW�(���3�P�E�e��u��E������E�d�    ËM�d�    Y__^[��]QËM�3��h��������M�3��Y���������U��� �EVWjY��s�}��E��E_�E�^��t� t�E� @��E�P�u��u��u������ ��U��3�@�} u3�]Ë�U��3�@�} u3�]Ë�U��3�@�} u3�]����������U��SVWUj j hh�u�4�  ]_^[��]ËL$�A   �   t2�D$�H�3����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�hpd�5    ��3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �ypu�Q�R9Qu�   �SQ�@��SQ�@��L$�K�C�kUQPXY]Y[� ��Ë�U��M�I�8 t@��u�I�E+�H]Ë�U�����3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5��3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w��d  ��;�t� ��  �P����Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5��SSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�d  ��;�th���  ���P���Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$�H��E�W�-���Y�u��$����E�Y�e�_^[�M�3�����Ë�U����u�M�����u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap��Ë�U��QQ��3ŉE�S3�VW�]�9]u�E� �@�E�5��3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w��b  ��;�t� ��  �P����Y;�t	� ��  ���؅�t��?Pj S������WS�u�uj�u�օ�t�uPS�u����E�S������E�Y�e�_^[�M�3��b���Ë�U����u�M��f���u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U���S�XBV���HD�M���u�����  �e� W�E�FPj1S�E�jP�T)�����FPj2S�E�jP�@)����FPj3S�E�jP�,)����FPj4S�E�jP�)����P��FPj5S�E�jP�)����FPj6S�E�jP��(��Vj7S��E�jP��(����F Pj*S�E�jP��(����P��F$Pj+Sj�E�P�(����F(Pj,S�E�jP�(����F,Pj-S�E�jP�(����F0Pj.S�E�jP�u(����P��F4Pj/S�E�jP�^(����FPj0S�E�jP�J(����F8PjDS�E�jP�6(����F<PjES�E�jP�"(����P��F@PjFS�E�jP�(����FDPjGS�E�jP��'����FHPjHS�E�jP��'����FLPjIS�E�jP��'����P��FPPjJS�E�jP�'����FTPjKS�E�jP�'����FXPjLS�E�jP�'����F\PjMS�E�jP�|'����P��F`PjNS�E�jP�e'����FdPjOS�E�jP�Q'����FhPj8S�E�jP�='����FlPj9S�E�jP�)'����P��FpPj:S�E�jP�'����FtPj;S�E�jP��&����FxPj<S�E�jP��&����F|Pj=S�E�jP��&����P����   Pj>S�E�jP�&������   Pj?S�E�jP�&������   Pj@S�E�jP�&������   PjAS�E�jP�w&����P����   PjBS�E�jP�]&������   PjCS�E�jP�F&������   Pj(S�E�jP�/&������   Pj)S�E�jP�&����P����   Pj�u��E�jP��%������   Pj �u��E�jP��%������   Ph  �u��E�jP��%������   Ph	  �u��E�j P�%����E���P���   ���   Pj1S�E�jP�%������   Pj2S�E�jP�q%������   Pj3S�E�jP�Z%������   Pj4S�E�jP�C%����P����   Pj5S�E�jP�)%������   Pj6S�E�jP�%������   Pj7S�E�jP��$������   Pj*S�E�jP��$����P����   Pj+S�E�jP��$������   Pj,S�E�jP�$������   Pj-S�E�jP�$������   Pj.S�E�jP�$����P����   Pj/S�E�jP�k$������   Pj0S�E�jP�T$������   PjDS�E�jP�=$������   PjES�E�jP�&$����P����   PjFS�E�jP�$������   PjGS�E�jP��#�����   PjHS�E�jP��#�����  PjIS�E�jP��#����P���  PjJS�E�jP�#�����  PjKS�E�jP�#�����  PjLS�E�jP�#�����  PjMS�E�jP�h#����P���  PjNS�E�jP�N#�����  PjOSj�E�P�7#�����   Pj8S�E�jP� #�����$  Pj9S�E�jP�	#����P���(  Pj:S�E�jP��"�����,  Pj;S�E�jP��"�����0  Pj<S�E�jP��"�����4  Pj=S�E�jP�"����P���8  Pj>S�E�jP�"�����<  Pj?S�E�jP�y"�����@  Pj@S�E�jP�b"�����D  PjAS�E�jP�K"����P���H  PjBS�E�jP�1"�����L  PjCS�E�jP�"�����P  Pj(S�E�jP�"�����T  Pj)Sj[�E�SP��!����P���X  Pj�u��E�SP��!�����\  Pj �u��E�SP�!����`  Vh  �u���E�SP�!����<�_^[�Ë�U��V�u���c  �v����v����v����v����v����v�y���6�r���v �j���v$�b���v(�Z���v,�R���v0�J���v4�B���v�:���v8�2���v<�*����@�v@����vD����vH����vL����vP�����vT�����vX�����v\�����v`�����vd�����vh�����vl�����vp����vt����vx����v|�����@���   ������   ������   ������   �x�����   �m�����   �b�����   �W�����   �L�����   �A�����   �6�����   �+�����   � �����   ������   �
�����   �������   ������@���   �������   �������   �������   �������   ������   ������   ������   ������   ������   ������   �x�����   �m�����   �b����   �W����  �L����  �A����@��  �3����  �(����  �����  �����  �����   ������$  ������(  ������,  ������0  ������4  ������8  �����<  �����@  �����D  �����H  �����@��L  �����P  �u����T  �j����X  �_����\  �T����`  �I����^]Ë�U��SV�u�~  W�X�tBhd  j�e&����YY��u3�@�I�Ƌ��R�����tW�G���W����YY��Ǉ�      ������   ;�t�   P�����   3�_^[]�2�8tSV�<0|<9,0�A8u�^[�<;u���X�@8u����U��V�u��tY�;X�tP�y��Y�F;\�tP�g��Y�F;`�tP�U��Y�F0;��tP�C��Y�v4;5��tV�1��Y^]Ë�U���SV�uW3��u��}�9~u9~u�}��}��X��e  jPj�8%����YY;�u3�@�  ���   jY��j���$��3�Y�E�;�u	S����Y�ыu�89~��   j�$��Y�E�;�u3�FS����u����YY���D  �8�v>SjV�E�jP�I�����CPjV�E�jP�5����CPjV�E�jP�!����C0PjV�E�jP�����P��C4PjV�E�jP�������tS�{���Y����k����C����0|��9��0�@�8 u��>��;u���N�F�> u���X���\��C�`��C����C0����}��C4�M��u3�@��M���t����   �=���tP�׋��   ��tP�ׅ�u���   �i�����   �^��YY�E����   �E����   ���   3�_^[��2�8tSV�<0|<9,0�A8u�^[�<;u���X�@8u����U��V�u����   �F;d�tP�� ��Y�F;h�tP�� ��Y�F;l�tP�� ��Y�F;p�tP� ��Y�F;t�tP� ��Y�F ;x�tP� ��Y�F$;|�tP� ��Y�F8;��tP�m ��Y�F<;��tP�[ ��Y�F@;��tP�I ��Y�FD;��tP�7 ��Y�FH;��tP�% ��Y�vL;5��tV� ��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}��X���  jPj�"����YY;�u3�@�  j�!��Y�E�;�u	S����Y���89~�4  j�!��Y�E�;�uS�����u�����Y�҉8�v8�CPjV�E�jP�@�����CPjV�E�jP�,����CPjV�E�jP�����CPjV�E�jP�����P��CPjV�E�jP������C PjPV�E�jP������C$PjQV�E�jP������C(PjV�E�j P�����P��C)PjVj �E�P�����C*PjTV�E�j P�����C+PjUV�E�j P�r����C,PjVV�E�j P�^����P��C-PjWV�E�j P�G����C.PjRV�E�j P�3����C/PjSV�E�j P�����C8PjV�E�jP�����P��C<PjV�E�jP������C@PjV�E�jP������CDPjV�E�jP������CHPjPV�E�jP�����P��CLPjQV�E�jP������t$S����S�����u������u�������������C����0|��9��0�@�8 u�� ��;u���N�F�> u���jY�X����E���   �	����   �I�u�K���   �I�K���   �I0�K0���   �@4�M��C43�@3��9}�t�M�����   ;�tP�����   ;�t#P����u���   ��������   �����YY�E����   �E����   ���   3�_^[���0���Hl;��t�P��Hpu��Q�����á�������ȋAl;��t�P��Qpu�Q�����   Ë�U���S�u�M������]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P��  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP������� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��=�� u�E����A#E]�j �u�u������]áD�øT�Ë�V���t��t;�tWj6Y���  P��M��Y_^Ë�U��V����Hpj Z���r�U���t0��t3��t��t�V-���    �R�������������Hp��P����^]á�����   ������   ������   �x��jhx��9(���u����   j��e��Y�e� �F��tP����u�F=0�tP�r���Y�E������[   �> t<j�e��Y�E�   �6�vM��Y���t�8 u=��tP��M��Y�E������&   �𭺉�FV����Y��'��Ëuj�id��YËuj�]d��YË�U��]�3���jh���l'���_����jj���YY���u��u�,���    3��[�O���HG���Gl��Gh�Fj��d��Y�e� �6�)L��Y�E������/   j��d��Y�E�   �v���E������   ���''��Ëu�j�c��YËu�j�c��Y��L���3�Ë�U��SW3�3�9]~"V�u���6�u�u�ci  ����uG;}|�^_[]�SSSSS�5P��̋�U��SVW�}h�   3�SW�w����u�����u3���   <.u1�F8t*jP���   jP���������u���   ��SSSSS��O��h(}V�]�Qi  ;��   �} �<0�u��@��   ��.t|PVj@�u�;�}u��@sh��_tcP�EVj@��@��}uQ��sL��t��,uCP�EVj��P�7�������u4��,�=������5����E�wh(}V�h  ��YY�k������_^[]�3�PPPPP�=�����U��SV�uV�u�u�]����3ۅ�uA�F@8tPh0}j�u�u�g��������   8^[tPh,}j�u�u�E�����]�SSSSS�N��̋�U���S3�ChU  �]��N��Y�E����=  W�x� ��vX�Q  h�l�5l|jSW������FX���E�l|�E�h4}SW�Vg  ������   �E��H�1�M��0����YY��t�e� �E��0�E�h�l�E��E��0jSW�������}��||��}� uU�FP����tP�Ӆ�u	�vP����Y�FT��tP�Ӆ�u	�vT�w���Y�E��fT �fL �FP�~H���Z3�PPPPP�M���u��M����FP�=�3�Y;�tP�ׅ�u	�vP�.���Y�FT;�tP�ׅ�u	�vT����Y�Fh�^T�^L�^P�^H_[�Ë�U���   ��3ŉE��ESV�uW�}��d����E��\�����`����N�����   ��T������   ���   K  ��X�����h�������  ��d��� ��  �} ��  �>CuS�~ uMh8}�u��d����c[������u'��tf�f�Gf�G��`�����t�  ��d����C  3�PPPPP�jL��V�`Z����   Y��P���;�s,V��h�������YY����   V��X�������YY����   ��L��� ��l���VP�����YY����   ��l���PSP�k  ������   �C��T������l���PW��h����������> t
��P���;�r��L�����l@PVW��X������������%���3�9�\���tjS��\����_�����9�`���tj��T�����`����A�������h����u��d����Z������u��h����VVVVV�����3��M�_^3�[�K����Ë�U����  ��3ŉE��ES��W��p�����h����;����S��\���P��P���Ph�   ��x���P��h�����������u3��M�_3�[�����������sH��x���P�P
��YY��u�CH�Ӎ�x���P�X����P��t����;��YY��l�����t��CH��p�����h����D���X���� ��H����Ak��jP��d�����8���P�����F��x���Q��t�����L�����l��������QP��X�������	  ��l�����X������CH��P����j��P���P��d�����������p����  ��\�����t��� �F���  ���  ��d������  �V;t6���t������d�����@����P�H��@�������t�����d���|��-��t�����t#����  ����  �P���  ���d����H��t���urj�v��x����vPjh�|jj ������� ��t<3���  f!�Ex���@��r�h�   �5����x���P�~  �����@���  ����   �F���  ���  ���   ��p���u	��\����F��p���k�V��h|Y��t1��h�����l����CH�+�����H���Y��X������L����F������h���T�t.��p�������4�����u�4�������sT������cL YY��p�����l�������    ���Y���3�PPPPP��G��̋�U���   ��3ŉE��ESV3ۋ�W��h���;�t;�tP����Y��  ɋD�H��  ǅp���   ��t���;���  �8L�0  �xC�&  �x_�  ��h<}W�0�  ��YY����   +ǉ�p�����   �;;��   ǅl���   �l|���p���PW�6��  ����u�6�U��Y9�p���t��l��������|~�Ch4}S�y`  ��3�YY;�u	�;;��   ��l���DWS��x���h�   P虾������uT��l�����h�����=x�����x���P�t���Y��t��t�����? t
G�? ����3�9�t�����   ��h����   VVVVV�YF��3��xSSSh�   ��x���QP�������;�t\�~H��t5�7��x���P����YY��t��x���P�������Y��u!�p������t���C����~�3�9�p���u9�t���t�3����M�_^3�[������Ë�U��}VWw$�} t3�GWj�����YY��u� ���    3�_^]�Wh�   ���YY���u	V�<���Y��Wh   �r��YY�F��u�6����V����Y�ً��������u�M��T���Y��u�6�A���6�A��V��������2�v��p�<��YY��t#�v������6��@���6�zA��V������3��
�F�8�F�8���>�����U��]� ���jhȨ����e� �}v����    �E��3��9  �������u��B���Np�e� 3�GWh�   �~��YY�؉]܅���   j�{X��Y�}��Nl�������e� �   �u�M���X���Y�E�����   �} thT��u����YY��t�=��j�%X��Y�E�   �~lSW��A��S��?�����Fpu?�P�u6�7h���A��YY������   ������   ������   �x��e� �   �.�]܋u�3�Gj�V��YËu�j�V��Y��S�i?��S��?��YY�E������   �E�����Ëu�fp�Ë�U����u�M������E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U��h  �u�	�  YY]Ë�U��h  �u��  YY]Ë�U��j�u���  YY]Ë�U��j�u�͏  YY]Ë�U��j�u躏  YY]Ë�U��j�u觏  YY]Ë�U��j�u蔏  YY]Ë�U��j�u聏  YY]Ë�U��h�   �u�k�  YY]Ë�U��h�   �u�U�  YY]Ë�U��j�u�B�  YY]Ë�U��j�u�/�  YY]Ë�U��j�u��  YY]Ë�U��j�u�	�  YY]Ë�U��h  �u��  YY]Ë�U��h  �u�ݎ  YY]Ë�U��hW  �u�ǎ  YY]Ë�U��hW  �u豎  YY]Ë�U��h  �u蛎  YY]Ë�U��h  �u腎  YY]Ë�U��j �u�r�  YY]Ë�U��j �u�_�  YY]Ë�U�츀   f9E���]Ë�U��h  �u�5�  YY��u	f�}_t]�3�@]Ë�U��h  �u��  YY��u	f�}_t]�3�@]Ë�U��h  �u��  YY��u	f�}_t]�3�@]Ë�U��h  �u�Í  YY��u	f�}_t]�3�@]Ë�U��UV�u�23�;�r;�s3�@�U�
^]Ë�U��E�jY#�U����  �yJ���B+ʃ����M�҅�t
3�]Ã<� u�@��|�3�@]Ë�U��ESVW�jY#�U����  �yJ���B�}+�3�B���3ۍ4;�r;�s3�C�4����t���Q3�;�r��s3�C��Hy�_^��[]Ë�U��QQ�e� SVW�}O�G�����G��%  �yH���@�ujY+�3�@���M�����   �������҅���<� u@��|��e�ǙjY#������  �yO���G�e 3�+�B����<;�r;�s�E   �M�<����t���Q3�;�r��s3�G����Hy��M��M������jY!�C;�}	+ˍ<�3��E�_^[�Ë�U��E�MjZ+�V�0�4��Ju�^]Ë�U��W�}3����_]Ë�U��3��M�<� u@��|�3�@]�3�]Ë�U��E�����UV����  �WyJ���B�e� �e �}��������E�    )U�S�֋M��#މ]������M]����]�M����E�}�]�|�jY��+Ѝ�[;�|�2�4���$� ��Iy�_^�Ë�U���<��3ŉE��E�M�M��H
�с� �  �MċH�M��H� S�]���  ���?  ��VW�U��M�E������u"3�3�9t��u@��|��  3��}𫫫�3  �e� �u��}䥥�¥�{�E�O�G�������W��  ��E�yJ���B�t��j3�Y+�@���M̅��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}܋99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U܉�M�yщMЋM̃����jY!�E�@;�}
�|��+�3��}� t�E��C�M���+S;�}3��}𫫫�  ;��  +Eԍu�}𥥋ș����4������  �yJ���B�e� �e� ��������E�    )U��ЋM��|����#ȉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���E�Y+�;�|��T����d�� ��Iy�{O�G�������W��  ��E�yJ���BjY+�3�B��M̅T����   �������օt����|�� uB��|��o�ǙjY#������  �yO���G�e� 3�+�B��L���9�4�u�;�r;�s�E�   �U܉�M����t�L����r3�;�r��s3�G�1��HyދEԋM̃����jY!T��@;�}
�|��+�3��K�A����4�Q����  �yJ���B�e� �e� ��������E�    )U��ЋM��|����#ȉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���E�Y+�;�|��T����d�� ��Iy�3�jX�N  ;�K��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�s33�@�   �su��e�������������с�  ��E�yJ���B�e� �e� ��������E�    )U��׋E��D����#ωMԋ���M�E؉D���EԋM����E��}��E�|ЋŰ�j���E�Y+�;�|�8�|����d�� ��Iy�3�jY+K�[��M���Ɂ�   ��u���@u�MȋU�q��
�� u�Mȉ1�M�_^3�[������Ë�U���8��3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=��O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�����+��;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5��N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��Ľ�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �Ľ;����   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�̽��3�@�   ̽�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+Ľ��M���Ɂ�   �ًȽ]���@u�M̋U�Y��
�� u�M̉�M�_3�[�}����Ë�U���8��3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=ؽO�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�Խ��+ؽ;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5ؽN�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��ܽ�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �ܽ;н��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy��н3�@�   ��e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+ܽ��M���Ɂ�   �ً�]���@u�M̋U�Y��
�� u�M̉�M�_3�[�,����Ë�U��� ��3ŉE��M�Q
�e� ��%�  �� �  V�q�E�Q�	��W�}�u��M���yd�����t\�J3�;�r��s3�F�e� �M�΅�t8�M�e� �L����r;�r��s�E�   �M�1�M�y҅�t
�E�   ���u��U���  f9M�u�E�   E�M��wf�G�E��_3�^�O����Ë�U��EV�0���W�x���0�4?�H������_�p�H^]Ë�U��E�P�HVW��������ΉH��������_�P�^]Ë�U���0��3ŉE��E3�S�]�S
V�MԉM��M�M��H
��3�� �  �u��  #�#֍4
W����  �u�f;���  f;���  ���  f;���  ��?  f;�w
3ɉH��  ����f��uF�uЅxu3�9Hu9uf�H
�  3�f;�uF�uЅ{u	9Ku9t��M�}��E�   �M�U�ɉU؅�~P���]܍�U����e� �ʋW��4
;�r;�s�E�   �}� �w�tf��m����M؃}� ��]�uЃ��E��M�}� ����  ���  f��~8�E�   �u*�M��]�U��e����ًM�������]�M�f���f��O�f��yH�����ɉM���E�t�EԋM��]�U��m�����ًM�������M�]�M�uσ}� tf�M�� �  f9M�w�U����� �� � u/�}��u&�e� �}��u�e� f9}�uf�M�F�f�E���E���E��  f;�sf�M�u�f��M�H�M��Hf�p
� 3�3�f9M���J��   ��� ���P��H�M�_^3�[�o����Ë�U���D��3ŉE��E�����`3҉M�9U��  }�]�����`�M�9Uu3�f�9U��  SVW�M�E�T�}��;��~  k�M܋ٹ �  f9r��}䥥��M�]��H
�UȉU��U�U��S
��3�� �  �uо�  #�#֍<
���}�f;��  f;���  ���  f;���  ��?  f;�w
3ɉH��  3�f;�u!G�@����}�u9pu90u3�f�H
��  f;�u#G�C����}�u9su93u�p�p�0�  �u̍u��E�   �M̋U�ɉUԅ�~S�SȉU��MċMċU���	�e� �ʋV��<
;�r;�s�E�   �}� �~�tf��E��m��Mԃ}� ��}؃��E��M��}� ����  f��~;�E�   �u-�u�M��e�������M����ʁ���  �u�M�f���f��M����  f��yB��������E�t�EȋM��]�U��m�����ًM������N�]�M�u�9u�tf�M�� �  f9M�w�U����� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�M�G�f�E���E���E��  f;�sf�M�}�f��M�H�M��Hf�x
� 3�3�f9M���J��   ��� ���P�H�3�9U�a���_^[�M�3��p����Ë�U���|��3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u����    �]'��3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$�WY�Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�q  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  �����`�E�;���  }�ع���E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^������ÍI ;S�S�S	TNT�T�T�T�T[UPU�T��U�����3ŉE��U�M�EV�uWR3�RRR�uQP�E�P��������E�VP�(�����(��u���M���_3�^�9����Ë�U��E�SVW�}��43�;�r;�s3�C�0��t�H�Q3�;�r��s3�F�P��t�@�H�W�43�;�r;�s3�C�p��t�@�OH_^[]Ë�U���t��3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uhX}�S3�PPPPP����3�f9U�t��   �u9Uu-hP}�;�u"9UuhH}�CjP�N-������u��C�h@}�CjP�1-������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع����`�ۉE�f�U�u�}�M���  ��y�����`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�����À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ������U��QQ�EV3��} 	 u:���u5��}��M���=  �=  f;�u95��t5�]��M�����  ���  t %����P�uV�n(������t
VVVVV�9��^�Ë�U��M3���tjX��t����t����t���� t����t   S��V�ʾ   #�W�   �   t!��   t��   t;�u��	��   #�t;�u   �   �E   _^[t   ]�3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   Ë�U��M3���?t2��tjX��t����t����t���� t����t   ]�3���yjXS�   VW��t����   t����   t����   t���   ��t   �ʾ `  #�t!��    t�� @  t;�u   ����_��@�  ��@^[t���  t��@u   �   �   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U��M3���?t2��tjX��t����t����t���� t����t   ]�h�  ��&  YË�U��QQV��}��E�3Ҿ   �?t)�tjZ�t���t���t��� t���tփ=�� tA�]��M�3���?t/��tjX��t����t����t���� t����t�����^�Ë�V�����0�������h�  �/&  Y��t�F�   t�`  �@$��  ^���%  3ɨ?t-�tjY�t���t���t��� t���t��   ��Ë�U��Q�]��e���U��M�3���?t2��tjX��t����t����t���� t����t   �Ë�U��QQ�e�]��M�3���yjXS�   VW��t����   t����   t����   t���   ��t   �ѿ `  #�t!��    t�� @  t;�u   ���ƾ@�  #΃�@t���  t��@u   �   �   �U�M#M��#��;���   �����P�E��$  Y�]��U�3���yjX��t����   t����   t����   t���   ��t   ��#�t$��    t�� @  t;�u   �	   ��#փ�@t���  t��@u   �   �   _^[�Ë�U��U��t<��}�E3ɨ?t-�tjY�t���t���t��� t���t��   �
V�u��t�����^]Ë�U��QQ�}���=�� ��   �E�3�V�   �?t)�tjZ�t���t���t��� t���t��]��e���U��M�3���?t/��tjX��t����t����t���� t����t��^�ÊM�3���?t2��tjX��t����t����t���� t����t   �Ë�U��E��SV3�W�   9U�V  ��}�f�]���tjZ��t����t����t���� t����t��   �ËȾ   #�t&��   t��   t;�u����   ���   #�t=   u��   ���   �é   t��   �]�E#E��#��;���   ��������E��m���}��U�3���tj[��t����t����t���� t����t��   �ʋ�#�t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �E��E�} ��  3�95���~  %�E��]�E��yj^�   t���   t���   t���   t���   t��   �ȿ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   �E���#E��#��;�u���   ����P�E�}   Y�]�M3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#˃�@t���  t��@u��   ���   ���   �M���E�0_3�^@[�Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ����������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95����  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��q  Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�Ë�U���SVW�}��������}f�]3���tjZ��t����t����t���� t����t��   �ˋ��   #�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   �é   t��   ���Ћ�#M#���E�;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U�3�95����  ���}��]�E��yj^�   t���   t���   t���   t���   t��   �ȿ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��V  Y�]��U�3���yjX��   t����   t����   t����   t���   ��t   ��#�t$��    t�� @  t;�u   �	   ��#Ӄ�@t���  t��@u   �   �   ��3M�E��� t   �_^[���������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��j
j �u��V  ��]Ë�U���uj
j �u��V  ��]Ë�U��]�������U��]�������U��j
j �u��Y  ��]Ë�U���uj
j �u��Y  ��]��������Q�L$+ȃ����Y�*Z  Q�L$+ȃ����Y�Z  ��U��QQ�EV�u�E��EWV�E��([  ���Y;�u����� 	   �ǋ��J�u�M�Q�u�P����E�;�u�����t	P����Y�ϋ������������D0� ��E��U�_^��jh ��s�������]܉]��E���u�/����  ����� 	   �Ë��   ��x;d�r�����  ������ 	   �B���ы����<�����������L1��t�P�Z  Y�e� ��D0t�u�u�u�u��������E܉U������� 	   �����  �]܉]��E������   �E܋U��������u��Z  YË�U���  �X  ��3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u�����8�����    �Y������  ������S����������L8$�����$�����?�����t��u'�M����u�����  �����    �����  �D8 tjj j V������V�>  Y����  ��D���  �����@l3�9H�� �����P��4�����3�;��`  ;�t8�?����P  �����4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P肾��Y��t:��4���+�M3�@;���  j��D���SP�]  �������  C��@����jS��D���P�`]  ������n  3�PPj�M�Qj��D���QP�� ���C��@����H������=  j ��,���PV�E�P��$���� �4������
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4�������  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����Z  Yf;�D����I  ��8�������� t)jXP��D����~Z  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4������C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4������i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �H���;���   j ��(���P��+�P��5����P��$���� �4�����t�(���;��������D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48�����t��(�����D��� ��8���������D�����8��� ul��D��� t-j^9�D���u������ 	   ������0�?��D��������Y�1��$���� �D@t��4����8u3��$�����    �����  ������8���+�0���[�M�_3�^�s�����jh ������]���u�Q����  �6���� 	   ����   ��x;d�r�*����  ����� 	   �e����ҋ����<����������D0��t�S��R  Y�e� ��D0t�u�uS�n������E������� 	   �����  �M���E������   �E�����Ë]S�S  YË�U�����h   � ���Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u�(���� 	   3�]Å�x;d�r����� 	   �c����ދȃ����������D��@]ø�á@�Vj^��u�   �;�}�ƣ@�jP����YY�����ujV�5@�����YY�����ujX^�3ҹ�������� ����p�|�j�^3ҹ �W������������������t;�t��u�1�� B��`�|�_3�^��X  �=�� t�3V  �5���¢��YË�U��V�u��;�r"��P�w��+�����Q�����N �  Y�
�� V���^]Ë�U��E��}��P�����E�H �  Y]ËE�� P���]Ë�U��E��;�r=P�w�`���+�����P���Y]Ã� P�|�]Ë�U��M�E��}�`�����Q�W��Y]Ã� P�|�]Ë�U��E��u�����    �t������]Ë@]�jh@��>���3�3�9u��;�u������    �@�������_�����j [�Pj�����YY�u�������P�QW  Y���EPV�u������P�{���E������PW��W  ���E������	   �E������������� Pj����YYË�U��EP�u�u�>X  ��]Ë�U��EP�u�u�BX  ��]Ë�U��EPj �u�*X  ��]Ë�U��EP�u�u�.X  ��]Ë�U��EPj �u�X  ��]Ë�U����U��3�9�������#щ��]á���3�9������Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v�h���j^�0�������V�u�M�肥���E�9X��   f�E��   f;�v6;�t;�vWSV�v���������� *   ����� 8]�t�M��ap�_^[��;�t&;�w �����j"^�0�I���8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p�H�;�t9]�j����M;�t��������z�P���;��s���;��k���WSV諔�����[�����U��j �u�u�u�u������]Ë�U����u�M���M��Q����E�P�u�E����   �E��uP�[�������u�E������}� t�M�ap��Ë�U��Q�M��j �u�  P�u�E�P��������u�E��Ã���Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�  �EPSj �u����M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U��j�u�u�u�u�u�u�������]Ë�U����ESV3ۋ���C�u��t�]tS�  Y����  �t�Etj�s  Y����x  ����   �E��   j�Q  �EY�   #�tT=   t7=   t;�ub��M����`���{L�H��M�����{,�`��2��M�����z�`����M�����z�P���P���������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�S  �M��]�� �����������}�E����M�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}����� "   ]������ !   ]Ë�U��3���p�;Mt
@��|�3�]Ë�t�]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���p�;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�  ����uV����Y�E�^�Ë�t��h��  �u(�  �u������E ���Ë�U��=X� u(�u�E���\$���\$�E�$�uj�/�����$]��J���h��  �u� !   �0  �EYY]Ë�U��QQ�=X� �E�E�]�u)�u�E����\$�E�\$�E�$�uj�������$�������h��  �u� !   ��  �E�YY�Ë�S��QQ�����U�k�l$���   ��3ŉE��s �CP�s�	�������u#�e��P�CP�CP�s�C �sP�E�P��������s�������=X� u+��t'�s �C���\$���\$�C�$�sP������$�P�~����$��  �s �  �CYY�M�3��&�����]��[Ë�S��QQ�����U�k�l$���   ��3ŉE��s(�C P�s�?�������u2�E��C����]����E�j �C P�CP�s�C(�sP�E�P��������s�5������=X� u,��t(�s(�C ���\$�C�\$�C�$�sP�6�����$�P�����$��  �s(�:   �C YY�M�3��L�����]��[�3�Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-\��]���t����-\��]�������t
�-h��]����t	�������؛�� t���]���Ë�U��Q�=�� t�]���e� �E���jh`�����3�9��tV�E@tH9t�t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%t� �e��U�E�������e��U�{���Ë�U��Q�=�� t�]��e���U���3�9��t�D�����?�3�9��t�1�����?����Ë�U��V3�95��t"�����M#M���E�����#��P����Y��^]Ë�U��������M��?�P�����Y]Ë�U���L��3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP葭��������  j覵��j��  W�E��۵��jW�E��е��jW�E��ŵ��jh  �E�趵����$�E�9]��  9]��v  ;��n  9]��e  9]��\  �Eԉ3��M܈@=   |�E�P�v�l����2  �}��(  �E�EЃ�~.8]�t)�E�:�t �x�����M�� �G;�~��8X�uڋE�SS�v   Ph   �u܉E�jS踂���� ����  �M��E�S�v��   W���   QW@Ph   �vS�X�����$����  �E�S�v�   WP�E�W@Ph   �vS�+�����$���b  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~U8]�tP�M�M�:�tD�I��҉M�;�(��H   ��M��E� �  f����M̋M��	9M�~�M���M�8Y�u�h�   ��   QP�ć��j��   PW赇���E�j��   QP裇�����   ��$;�tKP����u@���   -�   P�\������   ��   +�P�I������   +�P�;������   �0������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u�����Y���o�u��ܐ���u��Ԑ���u��̐���u��Đ��3ۃ�C�ˋ��   ;�tP�����   ���   ǆ�   uǆ�   �yǆ�    {ǆ�      3��M�_^3�[�ϋ���������ȋAl;��t�P��Qpu�������   Ë�U��E��u]������ ���   ]�袮���ȋAl;��t�P��Qpu�\����@��|����ȋAl;��t�P��Qpu�6����@��V����ȋAl;��t�P��Qpu�������3�Ë�U��MVW��t�}��u�����j^�0�6������A�U��u� ���> tFOu���t�+��B��tOu��u� ����j"Y����3�_^]��������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0�^I  YY��u
�M���9�yN�u��^;]~�_^3Ʌ���[��]ÁN  ����F�FË�U��Q��tP�> tKh�V�J���YY��t:h�V�9���YY��uj�E�Ph   �w�����t)�E���V����Y�E���j�E�Ph  �w�����u3��Ã}� u��p��Ë�U��3�f�Mf;���t����r�3�@]�3�]Ë�V3�� �A�B<w����
�A�<w�������t�Њ
��uڋ�^�3��
B��A|��Z~��a��w@��Ë�U���|��3ŉE�VW�}�����׋�������jx�E�P���   ���%���  PW�����u	!��   @�A�E�P���   ��G  YY��uW����Y��t���   ���   ���   ���   ���Ѓ��M�_3�^�E����� ��U��QV��j�E�P��%�  h      P�����u3��);u�t!�} t�E�0W�������V�������Y;�_t�3�@^�Ë�U���|��3ŉE�SVW�}�����׍��   ���������jx�E�P�F���%���  PW�Ӆ�u�f 3�@�c  �E�P�v�F  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6�F  YY��u�N  �~�R�FuO�F��t,P�E�P�6�G  ����u�6�N�~�����Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6��E  Y3�Y��u0�N   �F9^t
   �F�H9^t<�6�L���Y;Fu/Vj�9^u49^t/�E�P�6�E  YY��uVS������YY��t�N   9^u�~�F���Ѓ��M�_^3�[������ ��U���|��3ŉE�VW�}�����׍��   ������jx�E�P�F���%���  PW�����u!F@�\�E�P�6��D  YY��u
9Fu1Vj��~ u0�~ t*�E�P�6��D  YY��uVP���?���YY��t
�N�~�~�F���Ѓ��M�_3�^�Y����� �v�$�������Y�j@h1��F����Fu�f ��6������v�����@�F�����������f @�~ YY�FtjX�������jh3��F����F�   t�   t�u�f ��6���������@Y�FtjX������jh��F����Fu�f Ë�U��SVW蘧�����   �E��u�O  ��   ���@�_�t�8 tSjh8����������g ��t[�8 tV���t�8 t	�����������S���� ��   Wj@h0���������tf���t�; t	�������R�������I���t0�; t+S��������Y�j@h1��G����Gu�g ��G  ����G�G� ��   �u�ƃ����#��������u����   ����  ��   ����  ��   ��P�x�����   j�w�������   �E��tf�Of�f�Of�Hf�p�]��th�5���  f9u h�j@S��������t3�PPPPP����j@Sh  �w�օ�t,j@�C@Ph  �w�օ�tj
j��S�u�D  ��3�@�3�_^[]Å�t3Ʌ����D	��� �	+�t3Ʌ����D	��f�f;t1���+�t3҅��D���u�F�I+�t3Ʌ����D	��3�Ë;tg���+�t3҅��D���uP�F�Q+�t3҅��D���u5�F�Q+�t3҅��D���u�F�I+�t3Ʌ����D	��3�Ë�VW���N  �;tv���+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������t ����3�����  �A;Btw���B+�t3������D ����k  �q�B+�t3������D ����L  �q�B+�t3������D ����-  �q�B+�t3������t ����3����  �A;Btw���B+�t3������D �����  �q	�B	+�t3������D �����  �q
�B
+�t3������D �����  �q�B+�t3������t ����3����  �A;Btw���B+�t3������D ����Y  �q�B+�t3������D ����:  �q�B+�t3������D ����  �q�B+�t3������t ����3�����  �A;Btw���B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������t ����3����m  �A;Btw���B+�t3������D ����G  �q�B+�t3������D ����(  �q�B+�t3������D ����	  �q�B+�t3������t ����3�����  �A;Btw���B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������t ����3����[  �A;Btw���B+�t3������D ����5  �q�B+�t3������D ����  �q�B+�t3������D �����  �q�B+�t3������t ����3�����  �� �� �� �� ������׃���  �$���A�;B�tx�B��q�+�t3������D �����  �q��B�+�t3������D ����f  �q��B�+�t3������D ����G  �q��B�+�t3������t ����3����"  �A�;B�tw���B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������t ����3�����  �A�;B�tw���B�+�t3������D ����s  �q��B�+�t3������D ����T  �q��B�+�t3������D ����5  �q��B�+�t3������t ����3����  �A�;B�tw���B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������t ����3�����  �A�;B�tw���B�+�t3������D ����a  �q��B�+�t3������D ����B  �q��B�+�t3������D ����#  �q��B�+�t3������t ����3�����   �A�;B�tw���B�+�t3������D �����   �q��B�+�t3������D �����   �q��B�+�t3������D �����   �q��B�+�t3������t ����3���uy�A�;B�ti���B�+�t3������D ���uW�q��B�+�t3������D ���u<�q��B�+�t3������D ���u!�A��J�+�t3Ʌ����D	��3���u3�_^ËA�;B�tk���B�+�t3������D ���u��q��B�+�t3������D ���u��q��B�+�t3������D ���u��q��B�+�t3������t ����3���u��A�;B�tx�B��q�+�t3������D ����]����q��B�+�t3������D ����>����q��B�+�t3������D ��������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3����q����A�;B�tw���B�+�t3������D ����K����q��B�+�t3������D ����,����q��B�+�t3������D ��������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3����_����A�;B�tw���B�+�t3������D ����9����q��B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ����r����q��B�+�t3������t ����3����M����A��J�+��=���3Ʌ����D	��-����A�;B�tw���B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tx�B��q�+�t3������D ����}����q��B�+�t3������D ����^����q��B�+�t3������D ����?����q��B�+�t3������t ����3��������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ����k����q��B�+�t3������D ����L����q��B�+�t3������D ����-����q��B�+�t3������t ����3��������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3��������A�;B�tw���B�+�t3������D ����Y����q��B�+�t3������D ����:����q��B�+�t3������D ��������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3����m���f�A�f;B��]�����  �A�;B�tx�B��q�+�t3������D ����3����q��B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ����l����q��B�+�t3������t ����3����G����A�;B�tw���B�+�t3������D ����!����q��B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ����y����q��B�+�t3������D ����Z����q��B�+�t3������t ����3����5����A�;B�tw���B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ����g����q��B�+�t3������D ����H����q��B�+�t3������t ����3����#����A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������q��B�+�t3������D ����{����q��B�+�����3������D ������v�+��ޯ������U�z����̮���p�C�h�����ߡ~�^�1�V���Ԩ��̠{�K����U��VW�}�ǃ� ��  H��  H�l  H�!  H��  �M�ESj Z�2  �0;1tt�0�+�t3ۅ��Ít����+  �p�Y+�t3ۅ��Ít����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����e  �p�Y+�t3ۅ��Ít��3����B  �p;qtv�p�Y+�t3ۅ��Ít����  �p	�Y	+�t3ۅ��Ít�����  �p
�Y
+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����t  �p�Y+�t3ۅ��Ít����U  �p�Y+�t3ۅ��Ít��3����2  �p;qtv�Y�p+�t3ۅ��Ít����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����d  �p�Y+�t3ۅ��Ít����E  �p�Y+�t3ۅ��Ít��3����"  �p;qtv�p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít��3�����   �p;qtj�p�Y+�t3ۅ��Ít���uw�p�Y+�t3ۅ��Ít���u\�p�Y+�t3ۅ��Ít���uA�p�Y+�t3ۅ��Ít��3���u"��+�;�������σ���  �$�r����  �P�;Q�ti���Q�+�t3҅��t���u��p��Q�+�t3҅��t���u��p��Q�+�t3҅��t���u��p��Q�+�t3҅��t��3���u��P�;Q�tu���Q�+�t3҅��t����\����p��Q�+�t3҅��t����=����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����t����P�;Q�tu���Q�+�t3҅��t����N����p��Q�+�t3҅��t����/����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����e����P�;Q�tu���Q�+�t3҅��t����?����p��Q�+�t3҅��t���� ����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tm���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����D	��3���u3�[�  �P�;Q�tu���Q�+�t3҅��t����5����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t����p����p��Q�+�t3҅��t��3����M����P�;Q�tu���Q�+�t3҅��t����'����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t����b����p��Q�+�t3҅��t��3����?����P�;Q�tu���Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������p��Q�+�t3҅��t����r����p��Q�+�t3҅��t����S����p��Q�+�t3҅��t��3����0����P�;Q�tu���Q�+�t3҅��t����
����p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������I��@�+��8���3Ʌ����D	��(����P�;Q�tu���Q�+�t3҅��t����c����p��Q�+�t3҅��t����D����p��Q�+�t3҅��t����%����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����{����P�;Q�tu���Q�+�t3҅��t����U����p��Q�+�t3҅��t����6����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����m����P�;Q�tu���Q�+�t3҅��t����G����p��Q�+�t3҅��t����(����p��Q�+�t3҅��t����	����p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������Q��p�+�t3҅��t���������Q��p�+�t3҅��t���������Q��p�+�t3҅��t��3����^����P�;Q�tu���Q�+�t3҅��t����8����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3��������f�P�f;Q��f����Q��p�+�����3҅��T�����  ������P�;Q�tv�Q��p�+�t3҅��t����z����p��Q�+�t3҅��t����[����p��Q�+�t3҅��t����<����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t����l����p��Q�+�t3҅��t����M����p��Q�+�t3҅��t����.����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t����]����p��Q�+�t3҅��t����>����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����u����P�;Q�tu���Q�+�t3҅��t����O����p��Q�+�t3҅��t����0����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������p��Q�+�����3҅��T����������c����M�u��+�t3҅��D�����   �A�V+�t3҅��D�����   �A�V+�t3҅��D�����   �A�N+���   3Ʌ����D	��   �M�u��+�t3҅��D���ud�A�V+�t3҅��D���uI�A�N뤋M�u��+�t3҅��D���u �A�N�x����E�M� �	�g���3�_^]Ë�ɸ��U�>�N���ο��Ƿt�F�0�?��������f�8�!�1�߹������X�*��3�Ѹ������U��Q�e� S�]��u3��   V��ru�s���tn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9u�r��.�@��I��F�@��I��<�@��I��2�@��I��(�M�E�u�����t:u@FA;�r�3�^[��� �	+�����������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U��Q���  f9Eu3��ø   f9Es�E����A��E�Pj�EPj�����u!E��E��M#��Ë�U��]������U���u�u����YY]Ë�U����ES3�VW�E�N@  ��X�X9]�E  3ɉ]���}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�S3�;�r��s3�F�ډP��t
�U�B�U�P�M�U�E�} �X�P�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[�Ë�U���V�u�M���^���E�u��t�0��u$�~����    �԰���}� t�E�`p�3���  �} t�}|Ѓ}$ʃe� �M�S�W�~���   ~�E�P��jP�\���M������   ���B����t�G�ǀ�-u�M���+u�G�E���O  ���F  ��$�=  ��u*��0t	�E
   �6�<xt<Xt	�E   �#�E   �
��u��0u�<xt<Xu�_�����3��u���   �U����N�у�t�˃�0���  t0�K�����w�� ���;Ms�M9E�r(u;M�v!�M�} u#�EO�u �} t�}�e� �[�U��UщU��G늾����u�u=��t	�}�   �w	��u+9u�v&�މ���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�_[^�Ë�U��3�P�u�u�u9��uh���P������]Ë�U��j �u�u�u�u������]Ë�U��=�� j�u�u�uuh���j �f�����]Ë�U��j�u�u�u�u�I�����]Ë�U���<S�u�M��
\���M�E3�;�t�;�u%������    ����8]�t�Ẽ`p�3�3��O  9]t�}|Ѓ}$ʊV�u�W�]�]��M��x���   ~�E�P�E�jP�Y���uă���E����   �A��;�t��E�G�}�-�}�u�M��}�+u	�G�}��E�jY9]u%�}�0t	�E
   �7�<xt<Xt	�E   �$�M9Mu�}�0u�<xt<Xu�G���E��}��E�R��Wj�j��U�迦���]����   �M܉E�U�M����C�Ѓ�t���0�%  tP�A�<��w�� �p�;us;�M��M;M�rQw�E�;E�rG�E�9E�u;M�u3�;E�r3w;u�v,�M�} u;�E�M��uA3�9Et�M�M��E�E��   Q�u��u�W�N  3��щE�U��E�� �E��E��E��������   ��u'�uT��t9]�wr�}� w��u>9u�r9w�}��v1跆���E� "   t
�M���M����Et	�e� �]���M���u��E_^��t�M���Et�E�M��؃� �ىE�M��}� t�Ẽ`p��E�U�[�Ë�U��3�P�u�u�u9��uh���P�=�����]Ë�U��j �u�u�u�u� �����]Ë�U��=�� j�u�u�uuh���j �������]Ë�U��j�u�u�u�u�������]���������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��EVW��xY;d�sQ���������<�������<�u5�= �S�]u�� tHtHuSj��Sj��Sj������3�[������ 	   � ����  ���_^]Ë�U��MS3�VW;�|[;d�sS��������<�������D0t6�<0�t0�= �u+�tItIuSj��Sj��Sj�������3��蒄��� 	   蚄������_^[]Ë�U��E���u�~����  �c���� 	   ���]Å�x;d�r�Z����  �?���� 	   蕩���Ջ������������Dt͋]�jh���I���}����������4����E�   3�9^u5j
����Y�]�9^uh�  �FP�0���u�]��F�E������0   9]�t�������������D8P����E��
���3ۋ}j
萻��YË�U��E�ȃ����������DP�|�]�jh���~���M��3��}�j�z���Y��u����a  j�(���Y�}��}؃�@�;  �4�������   �u�����   ;���   �Fu[�~ u8j
�߻��Y3�C�]��~ uh�  �FP�0���u�]���F�e� �(   �}� u�^S����FtS�|���@냋}؋u�j
莺��YÃ}� u��F��+4�����������u�}��uyG�,���j@j �4r��YY�E���ta������d� ���   ;�s�@ ���@
�` ��@�E������}�����σ��������DW�����Y��u�M���E������	   �E��E}���j�й��Y�jhȩ��|��3��}�2��Et�� �E @  t�ˀ�E�t���u�4�;�u���P葁��Y�����|��Ã�u��@���u����������u���u�;����    �C����8�}��uV����YY�����������ƃ�����\��T$�"��	�D$� �E�   �E������   9}��i������e����u3�9}�u�����΃��������D� �V�,���YË�U��Q�=���u�   ������u���  ��j �M�Qj�MQP�����t�f�E��jh��{��j�T���Y�e� �u����Y���E��E������
   f�E��{���j�2���YË�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��S���E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P�Fa��YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p������E�u�M;��   r 8^t���   8]��f����M��ap��Z����B��� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p������:���뺋�U��j �u�u�u�������]�jh��z��3ۉ]�j�ٷ��Y�]�j_�}�;=@�}T�����9�tE���@�tP�  Y���t�E��|(������� P�<�����4��(L��Y�����G��E������	   �E���y���j�f���YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV����YP蹦����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV����P�4  Y��Y��3�^]�jh(���x��3��}�}�j芶��Y�}�3��u�;5@���   �����98t^� �@�tVPV脨��YY3�B�U�������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u����4�V荨��YY��E������   �}�E�t�E��Qx���j�ܴ��Y�jhP���w��3�9uu	V����Y�'�u萧��Y�u��u����Y�E��E������	   �E���w����u�֧��Y�j�����YË�U��V�uV�'���P����YY��t|�a����� ;�u3���Q�����@;�u`3�@����F  uNSW�<����? �   u S�k��Y���u�Fj�F�X�F�F��?�~�>�^�^�N  3�_@[�3�^]Ë�U��} t'V�u�F   tV�`����f�����f �& �f Y^]�jhp���v��蠥���p �u�3�9E����u�m{���    �à������<V�J���Y�e� V��������u�u�uV�U�E�VW�j������E������   �E��v��Ëu�V�x���YË�U���u�u�uh���c�����]Ë�U���u�u�uh��F�����]Ë�U���u�u�uhN��)�����]Ë�U���uj �uh��������]Ë�U���uj �uh��������]Ë�U���uj �uhN��������]Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U���E��%�  -�  �]Ë�U���E�E�M��%�  �����PQQ�$������]Ë�U��QQ�M�E�E�]������  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$�m������&Q���EQQ�$�X����U�����  �����  �E�]Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M��K���]��u#�Gx���    蝝��8]�t�E��`p������V�u��u$�x���    �r����}� t�E��`p������R�E��x uVS�M���YY�1+�W�3�M�QP�̣������M�QP轣����F��t;�t�+���_�}� t�M��ap�^[�Ë�U��3�9��u'9Eu�w���    ��������]�9Et�]�����P�u�u�������]Ë�U����} SVW��   �u�M��sJ���]��u'�4w���    芜���}� t�E��`p������   �u��tҿ���9}v!��v���    �R����}� t�E��`p����]�E��x u�uVS�N'  ���}� tA�M��ap��8+��3�M�QP蟢������M�QP萢����F�Mt��t;�t�+����3�_^[�Ë�U��3�9��u09Eu�ev���    軛������]�9Et�}���w�]��&  P�u�u�u�������]Ë�U��SV��3�;�u�v��j^�0�n������   W9]w��u��j^�0�R������u3�9]���A9Mw	��u��j"�ۋM�����"wɋ�9]t3�C�-�N�؋�3��u��	v��W���0�AC��t;]r�;]r� �� I���I�G;�r�3�_^[]� ��U��}
�Eu
��yjj
�j �u�u�M����]Ë�U��3��}
u9E}@�MP�u�E�u�����]Ë�U��M�Ej �u�u�����]Ë�U���3�V;�u��t��j^�0�I�������   9Mv�3�9M���@9Ew	��t��j"�ӋE�����"w��ES�]�M���9Mt����-�w�E�   �؉u�M�u�uPS肓���]��؋�	v��W���0��M�FA�M���u��t;MrȋM�[;Mr� �Et��j"Y����L���� N�E���N�@�E;�r�3�^�� ��U��3��}
u9E
|9Es3�@W�}P�u�u�u�u�����_]Ë�U��W�}j �u�u�u�u�����_]�������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� 3�PPjPjh   @h �������á�����t���tP���Ë�U��V�uW�����u�?s���    蕘����D�F�t8V�����V���^%  V����P�$  ����y�����F��tP�@���f Y�f ��_^]�jh���n���M��3��u������u��r���    ���������F@t�f �E��)n���V菝��Y�e� V�<���Y�E��E������   �ԋuV�ܝ��Y�jh���m���]���u�[r��� 	   ����   ��x;d�r�<r��� 	   蒗���ڋ����<����������D��t�S�����Y�e� ��Dt1S�x���YP�����u����E���e� �}� t��q���M���q��� 	   �M���E������   �E��-m��Ë]S�(���Y��A@t�y t$�Ix��������QP����YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U��Q�C@V����E�t�{ u�E�>�' �} ~0�E� �M���n����E�>�u�?*u�˰?�X����} Ճ? u�E��^�Ë�U���  ��3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������C���tp����������u+�ep���    軕�������� t
�������`p�����a  �F@u^V����Y�@����t���t�ȃ��������������A$u����t���t�ȃ������������@$��q���3�;��g��������������������������������������
  C������9�������
  �B�<Xw��������3�������k�	��0�j��^������;������jY;�� 
  �$�3�3����������������������������������������������	  �� tH��t4+�t$HHt����	  	������	  �������	  �������	  �������   �	  �������	  ��*u,�������������������l	  �������������Z	  ������k�
�ʍDЉ������?	  ������ �3	  ��*u&�������������������	  ��������	  ������k�
�ʍDЉ�������  ��ItU��htD��lt��w��  ������   ��  �;luC������   �������  �������  ������ �  �<6u�{4u�������� �  �������o  <3u�{2u������������������M  <d�E  <i�=  <o�5  <u�-  <x�%  <X�  ������ ������ ������P��P��N��Y��������Yt"�������������u����C��������������������������S����  ��d��  �U  ��S��   tL��AtHHt$HHtHH��  �� ǅ����   �������S  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ��u�Լ������������ǅ����   ��  ��X�  HHt+���  HH��  ��������������  ������t0�G�Ph   ������P������P�m�������tǅ����   ��G�������ǅ����   �������������y  �����������t<�H��t5������   � ������t�+���ǅ����   �4  ������ �(  �м������P����Y�  ��p�6  �"  ��e��  ��g��   ��itx��nt*��o��  �������������������tl������   �`�������������p���������J��������� tf������f���������ǅ����   �>  ������������@ǅ����
   �������� �  ��  ��G��W��	  ������������@������ �������   ������������}ǅ����   �ju��gucǅ����   �W9�����~�������������   ~=��������]  V�Y��������Y��������t���������������
ǅ�����   ��5�����������G�������������P��������������������P������������SP�5 ����Ћ���������   t������ u������PS�5,�����YY������gu��u������PS�5(�����YY�;-u������   C������S������������������*��s�t���HH�[�������  ������ǅ����'   �������ǅ����   �5���������Qƅ����0������ǅ����   ������   �������� t��������@t�G���G����G���@t��3҉�������@t��|��s�؃� �ځ�����   ������ �  ����u3������� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPWS讆����0�������؋���9~������N뽍E�+�F������   ������������tc��t�΀90tX�������������0@�@If�8 t����u�+��������(��u�м�������������I�8 t@��u�+����������������� ��  ��������@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����+�������������u%���������������� O������������t���������������������������P����������������YYt.������u%��������������˰0O�����������t��ヽ���� ������tu��~q�������������������Pj�E�P������P��蓔������u69�����t.�������������������E�P�������s��������� YYu��#��������������P�������������E���YY������ |2������t)�������������������� O�����������t��߃����� t��������2�������� Y���������������t������3����d��������� t����������������� t
�������`p��������M�_^3�[��-���ÍI ������F����������U��S�]V�u�F<p�  ��p��   <st<St3��3�B��st	��St3��3�A����   ����   �d:�tM<it-<ot)<ut%<xt!<Xt:�t��it��ot��ut
��xt��Xu^:�t<it<ot<ut<xt<Xt3��3�A:�t��it��ot��ut��xt	��Xt3��3�@;�uK�F��3M��   u;3E� u4�3�;M���5;�u$�N�U�  #����#��������;�u3�@�3��	3�:�����^[]��A@t�y t$�Ix��������QP����YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U��Q�C@V����E�t�{ u�E�>�' �} ~0�E� �M���n����E�>�u�?*u�˰?�X����} Ճ? u�E��^�Ë�U��E� ��A��Q�]Ë�U����  ��3ŉE��ES�]V�uW�u3���������d�����������H�����������`�����L�����X����5�����������h����Db����D���;�u+�5b���    苇�������� t
�������`p�����R  �F@u^V�ԍ��Y�@����t���t�ȃ��������������A$u����t���t�ȃ������������@$��q���;��i�����������(���������������u9�������  3���(�����l��������������������x������T�����P�����p������������������E  ���������G������ ��|�����  �C�<Xw�������3��3�3���T���k�	��0�3���F��T���;���   �?%��   �������uQj
��h���PW�5�������~2��h����8$u'������ uh@  ������j P��#����������������� 3�9�����u]j
��h���PW�������h�����H������ �Q��������|���u(��������9$�������d�����;�l���~��l�����3ҋ�T����$�R����������r  ��9�����u9������\  9�������  ���������  �>  ���������8�����L�����p�����`�����������X����  �Ã� tI��t5��t%HHt����  ��������  ��������  	�������  �������   �  �������  ��*��   9�����u�������������@��   j
��h���PW�y�����h�����H������ �Q��|���uL��������9$�����������d�����;�l���~��l������Ŵ����9 ��   ������j*V�3  ���Ÿ���� 3҉�p���;���  ��������p�����  ��p���k�
�ˍDЉ�p�����  ��������  ��*��   9�����u�������������@��<j
��h���PW������h�����H������ �Q��|����������Ÿ���� 3҉�����;��T  ��������H  �1Ƅż���*��������������,  ������k�
�ˍDЉ������  ��ItU��htD��lt��w��  ������   ��  �?luG������   ��|�����  ��������  ������ �  �<6u�4u�������� �  ��|����  <3u�2u�������������|����q  <dt{<itw<ots<uto<xtk<Xtg��T�����X��� ������P��P�P>��YY��t,��d����������������G��������|������K����؋�d������������������  ������   ��  �Ã�d��  ��  ��S��   tA��AtHHt HHtHH��	  �� ��8����������i  ������0  uz������   �n������0  u
������   ���������u����9�������  �������������@���  ��X��  HH�K  ����  HH�%	  3�F3ҋ�������  ��   9�����u�������������@��f��������c�����9�����uC��Ŵ���9u�   ��ż�����������  W������jQ�k�������������  ��Ÿ���� Ph   ������P��x���P蒉������tq��L����i9�����u�������������@��B��������c�q����9�����u��Ŵ���9u�1�V���W������V�e�����Ÿ���� ��������x�����������������  9�����u�������������@��&��������c������9������  ��Ÿ���� ;�tV�H;�tO������   � ������t/�+�����X����u  �   ��������ż�����������\  ��X����K  �м������P行��Y�4  ��p��  ��  ��e�"  ��g��   ��i��   ��nt3��o�  ������3�Fǅ\���   ��y��   ������3��  3�9�����u�������������p��&��������c������9�������  ��Ÿ����0�D���������������� tf������f���������ǅL���   �]  3�F3҃�����@ǅ\���
   �f  3�F3҃�����@9�����uZ9�����uR��������c�M������Ŵ���9u�   ��ż�������������������jQ��������������  �������   ��������@���9�����}ǅ����   �gu������guZ�������T9�����~��������   9�����~7��������]  V�G��3�Y��P�����t��������@������
�������3�9�����u����������������@���,����'������c�G������������Ÿ������,����@�5����0���������P��8���������������P��@�����,���SP�5 ����Ћ���������   t������ u������PS�5,�����YY������gu��u������PS�5(�����YY�;-u������   C������S����ǅ����   ǅH���   �)��s�����HH��������  3�FǅH���'   3��������ǅ\���   t��H���Qƅt���0��u���ǅ`���   �������� �  tv9�����u��������Q����������  ��������c�����9�������   ���Ŵ���9u�   ��������ż�����������f  S������j������   t[9�����t���������c�o���9�����u#���Ŵ���9u�   �S������j�a������������Ÿ�����Q�:  �� ��   ��@tM9�����u�������������@���   ��������c�����9�����tJ���Ÿ���� �   �1����9�����u�������������@����������c�����9�����u���Ŵ���9t�S�7������������Ÿ���� �A��@t?9�����u�������������@��"��������c�I���9�����t����Ÿ���� ��B9�����u�������������@��&��������c�
���9������`������Ÿ���� 3���@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!�`��������������������������t-��\����RPSW�r����0��@������ڃ�9~�H����N뽍�����+�F������   ��x�����������   ��t�΀90��   �������������0@�   ��������c������9�����u"��Ŵ���9����������������j�������Ÿ���� ������  ������t4;�u�Լ��������������X����	If9t��;�u�+��������,9�����u�м�������������I�8 t@;�u�+�������x���������u������ ��  ��L��� ��  ��������@t5��   t	ƅt���-���t	ƅt���+���tƅt��� ǅ`���   ��p���+�x���+�`�����@�����u%�����d���������� O�W����������t�����`�����D�����d�����t���P����������������YYt.������u%��@�����������˰0O������������t��ヽX��� ��x���tu��~q��������\������\���Pj�E�P��4���P����������u69�4���t.��4�����D�����d����E�P�������������\��� YYu��#����������D���P����������������YY������ |2������t)��@������d���������� O�!����������t��߃�P��� t��P����4����P��� Y��|�������������6���3�9�T���t��T�������������uW9�����uO9�l���|G�������������H�ItItItItItItII������������F��������;�l���~�������������}3��E��������� t
�������`p��������M�_^3�[�����Ð�H�x�������u�����������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV����Y���tP�����u	���   u��u�@Dtj�f���j���]���YY;�tV�Q���YP�����u
������3�V����������������Y�D0 ��tW�N��Y����3�_^]�jhЪ�I���]���u�|N���  �aN��� 	   ����   ��x;d�r�UN���  �:N��� 	   �s���ҋ����<����������D0��t�S�����Y�e� ��D0tS�����Y�E����M��� 	   �M���E������   �E��PI��Ë]S�K���YË�U��V�u�F��t�t�v�U���f����3�Y��F�F^]��%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���% ��%��%��%��%��%��%��%��% ��%$��%(��%,��%0��%4��%8��%<��%@��%D��%H��%L��%P��%T��%X��%\��%`��%d��%h��%l��%p��%t��%x��%|��%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%���%�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̍M��H����|����|����,����q��������f����<����[����d����P����L����E���M��=���M��5���T$�B�����3��������"���M������T$�B�J�3��h���T���"���M������M��E���M��M���M�����M�����M�����M������M������M�m����M�����T$�B��X���3������x��R"���M��?���T$�B�J�3���������/"�����̋M��x���M���m���T$�B�J�3�����(���!���̋M��H���T$�B�J�3�����T���!��������������̍M�����M������T$�B�J�3��H������!���T$�B�J�3��-�����!��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������h�#�N��Y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̃=�� uK�����t����Q<P�B�Ѓ����    �����tV����+��V�
V�������    ^��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                          p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        [!51u!                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��                                                                                                                                                                                                                                                                �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                /��T       X   � {                                                                                                                                                                 	              	            	              	         ?             @                  �   &   ��������5            4  �������5            4  �������                e:\cinema4d\cinema4dr13\resource\_lib_welter\include\mycontainersmem.h                  p��  � P� P ` p � � � � � � � �� �� �� �� �� Ѐ ��  �  �                     e:\cinema4d\cinema4dr13\resource\_lib_welter\include\dynamicarray.hpp                         �?        e:\cinema4d\cinema4dr13\resource\_lib_welter\include\mycontainersarray.h                �'  � P�  � � p �� �� � � � � �� �� �� ��  � Ѐ P�  �  � �                        e:\cinema4d\cinema4dr13\plugins\pointcollapse\source\pointcoll.cpp              l�  � P� p � p P B � � O b � �� �� �� ��  � Ѐ P�  �  � .                     toolpointcollapse       pcoll.tif         �?    e:\cinema4d\cinema4dr13\resource\_api\c4d_resource.cpp  #   M_EDITOR    Е�~ res ����MbP?��,� �  � t� � e:\cinema4d\cinema4dr13\resource\_api\c4d_baseobject.cpp    ���� ��� X� �       �?e:\cinema4d\cinema4dr13\resource\_api\c4d_general.h %s  e:\cinema4d\cinema4dr13\resource\_api\c4d_general.cpp   %s(%d): %s     e:\cinema4d\cinema4dr13\resource\_api\c4d_file.cpp  e:\cinema4d\cinema4dr13\resource\_api\c4d_basebitmap.cpp    �������������e:\cinema4d\cinema4dr13\resource\_api\c4d_libs\lib_ngon.cpp e:\cinema4d\cinema4dr13\resource\_api\c4d_string.cpp     B   KB  MB       P? GB e:\cinema4d\cinema4dr13\resource\_api\c4d_pmain.cpp �� �e:\cinema4d\cinema4dr13\resource\_api\c4d_gv\ge_mtools.cpp  �P�4�������        �0w,a�Q	��m��jp5�c飕d�2�����y�����җ+L�	�|�~-����d�� �jHq���A��}�����mQ���ǅӃV�l��kdz�b���e�O\�lcc=���� n;^iL�A`�rqg���<G�K���k�
����5l��B�ɻ�@����l�2u\�E���Y=ѫ�0�&: �Q�Q��aп���!#ĳV���������(�_���$���|o/LhX�a�=-f��A�vq�� Ҙ*��q���俟3Ը��x4� ��	���j-=m�ld�\c��Qkkbal�0e�N b��l{����W���ٰeP�긾�|�����bI-��|ӌeL��Xa�M�Q�:t ���0��A��Jו�=m�Ѥ����j�iC��n4F�g�и`�s-D�3_L
��|�<qP�A'�� �%�hW��o 	�f���a���^���)"�а����=�Y��.;\���l�� �������ұt9G��wҝ&���sc�;d�>jm�Zjz���	�'� 
��}D��ң�h���i]Wb��ge�q6l�knv���+ӉZz��J�go߹��ﾎC��Վ�`���~�ѡ���8R��O�g��gW����?K6�H�+�L
��J6`zA��`�U�g��n1y�iF��a��f���o%6�hR�w�G��"/&U�;��(���Z�+j�\����1�е���,��[��d�&�c윣ju
�m�	�?6�grW �J��z��+�{8���Ғ�����|!����ӆB������hn�����[&���w�owG��Z�pj��;f\��e�i�b���kaE�lx�
����T�N³9a&g��`�MGiI�wn>JjѮ�Z��f�@�;�7S���Ş��ϲG���0򽽊º�0��S���$6к���)W�T�g�#.zf��Ja�h]�+o*7������Z��-   ��ư>      @      @{�G�z�?:�0�yE>e:\cinema4d\cinema4dr13\resource\_lib_welter\source\uvcomponentsmesh.cpp            �9��    �9�Cinner vertices  selected vertices   neighbored vertices border vertices -comp         Y@+ȘU                    e+000   r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
         R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            �`   �`	   H`
    `   �_   H_    _   �^   8^   �]   x]   ]   �\   x\   �[    H[!   XYx   4Yy   Yz   �X�   �X�   �XM i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     @���K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �             ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �        ]�[W
bad exception   H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun  Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    \mTmHm<m0m$mmmm�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l|lxltlplllhldl`l\lXlTlPlLlHlDl@l<l0l$lll�k�k�k�k�kxkXk8kk�j�j�j�jpj`j\jTjDj jjj�i�i�i�ipiHii i�h�h�h`hDh�l0hh h�g�g�����ĖȖ	��6�|���
�3�^�z�לۜ� ??     {flat}  {for    `non-type-template-parameter    unsigned    long    int     short   char    void    <ellipsis>  ... ,<ellipsis> ,...     throw( )[  s   '   `template-parameter NULL    cli::pin_ptr<   cli::array< void    ''  `anonymous namespace'   `   generic-type-   template-parameter- ::  `unknown ecsu'  union   struct  class   enum    coclass     cointerface     )   extern "C"  [thunk]:    public:     protected:  private:    virtual     static  `template static data member destructor helper' `template static data member constructor helper'    `local static destructor helper'    `adjustor{  `vtordisp{  `vtordispex{        }'  }'  const   volatile    CV:     volatile     volatile   const   signed  double  bool    <unknown>   wchar_t UNKNOWN __int128    __int32 __int64 __int16 __w64   __int8  float   long    int short   char    std::nullptr_t  GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L     SystemFunction036   A D V A P I 3 2 . D L L     ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          ���W
Unknown exception   ���W
�3W
<�wW
csm�               �                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  X|    |)L|T��@|T���4|T��"(|T�� |T�o	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., .   _   ;   C   =;  1#QNAN  1#INF   1#IND   1#SNAN  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   modf    fabs    floor   ceil    tan cos sin sqrt    atan2   atan    acos    asin    tanh    cosh    sinh    log10   log pow exp united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    $�ENU �ENU ��ENU ��ENA �NLB ܂ENC ؂ZHH ԂZHI ̂CHS ��ZHH ��CHS ��ZHI |�CHT l�NLB X�ENU L�ENA <�ENL 0�ENC �ENB �ENI  �ENJ �ENZ ܁ENS ��ENT ��ENG ��ENU ��ENU ��FRB |�FRC h�FRL X�FRS H�DEA 4�DEC  �DEL �DES  �ENI ��ITS �NOR ЀNOR ��NON ��PTB ��ESS ��ESB p�ESL \�ESO H�ESC ,�ESD �ESF �ESE �ESG �ESH �ESM �ESN �ESI �ESA �ESZ xESR dESU TESY @ESV 0SVF (DES $ENG  ENU ENU USA GBR CHN �~CZE �~GBR �~GBR �~NLD �~HKG �~NZL �~NZL �~CHN �~CHN �~PRI �~SVK �~ZAF x~KOR h~ZAF \~KOR H~TTO $GBR 8~GBR (~USA  USA 6-OCP ACP Norwegian-Nynorsk   C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               RSDS�I3����B��D���	   E:\Cinema4D\cinema4dr13\plugins\PointCollapse\pointcollapse.pdb                                                                                                                                                                                                                                                                                                  ���               ��    ��̔     �       ����    @   ��        �        ����    @   �                   �    ̔                8�$�               8�    H���̔    8�       ����    @   $�                    `���               ��    ��H���̔    `�       ����    @   ��                    ��            ����           ��    ��        ����    @   ��            ��@�           P�X�    ��        ����    @   @�            ����           �����    ��       ����    @   ��            ذԖ           ���    ذ       ����    @   Ԗ             � �           0�<��     �       ����    @    �            $�l�           |����    $�       ����    @   l�            H���           ȗЗ    H�        ����    @   ��            d� �           ��    d�        ����    @    �            ��H�           X�d��    ��       ����    @   H�            ����           ����    ��        ����    @   ��            бܘ           ���    б        ����    @   ܘ            �$�           4�@�\�    �       ����    @   $��        ����    @   x�           ��\�                �x�            ؼ��           șԙ\�    ؼ       ����    @   ��            ���           � �\�    ��       ����    @   �            �P�           `�p� �\�    �       ����    @   P�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    % & �P �� p z �  1 c � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "�	   �                       ����     (   3   >   I    T    _    j    r�����"�   L�                       "�
   ��                       �����    �   �   �   �   �    �   �   �   ����)"�   �                       ����P    X"�   �                       �����"�   L�                       �����    �"�   x�                           ����    ����    ����    �    ����    ����    ����_ p     ����    ����    ����    �!    ����    ����    ����    �6    ����    ����    ����    �7    ����    ����    ����    �7    ����    ����    ����    29    ����    ����    ����    �9    ����    ����    ����    �@����    �@����    ����    ����    iB����    uB����    ����    ����    �H    ����    ����    ����    �\    h\r\����    ����    ����N]W]    ����    ����    �����_`    ����    ����    ����.`8`    ����    ����    ����``j`    ����    ����    �����`�`@           \a����    ����                  �"�   ��   �                   ����    ����    ����    Lc    �b�b����    ����    ����3e7e    ����    ����    �����e�e    
[    ��   ��ܦ    �    ����       l    �    ����       �����    ����    ����4m8m    ����    ����    �����m�m    ����    ����    ����    �p    ����    ����    ����    �t    ����    ����    ����    |x    ����    ����    ����     �    ����    |���    ����    ��    ����    |���    ����    B�    ����    ����    ����    ��    ����    ����    ����    t�    ����    ����    ����    �    ����    ����    ��������    ����    ����    ����    �(����    �(����    ����    ����    _)����    k)����    ����    ����    �6        O6        a6    ����    ����    ����    �v    ����    ����    ����    q~    ����    ����    ����    ��    ����    ����    ����ƍ�    ����    ����    ����    |�    ����    ����    ����    A�        }�����    ����    ����    3�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    5�        �����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    Y�    ����    ����    ����    6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        /��T    �          � � � � �   pointcollapse.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �X    .?AVToolData@@      �X    .?AVBaseData@@      �X    .?AVDescriptionToolData@@       �X    .?AVPcToolData@@        �X    .?AVGeSortAndSearch@@   �X    .?AVNeighbor@@  �X    .?AVDisjointNgonMesh@@  �X    .?AVTranslationMapNewSearch@@   �X    .?AVTranslationMapSearchN@@ �X    .?AVTranslationMapSearch@@  �X    .?AVGeToolNode2D@@  �X    .?AVGeToolDynArray@@    �X    .?AVGeToolDynArraySort@@    �X    .?AVGeToolList2D@@  u�  s�      �X    .?AVtype_info@@         N�@���D        sqrt    ����������   ��������    �����
                                                                                           	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 �X    .?AVbad_exception@std@@ �X    .?AVexception@std@@                                                                                                                                                                                                                                                                                                                                         abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     0��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����C   �g�g�g�g�g�g�g�g�g�g�gxgpgdg`g\gXgTgPgLgHgDg@g<g8g4g,g gggPgg g�f�f�f�f�f�f�f�f�f�f	         �f�f�fxfpfhf`fPf@f0fff�e�e�e�e�e�e�e�e�e�e�e�e�e�ete`eTeHe�e<e0e ee�d�d�d�d�d�d�dtd                                                                                           T�            T�            T�            T�            T�                              X�        u�y {X�����0�                                                                                                                                                                                                                                                                                              Ps@s�X    .?AVbad_cast@std@@  �X    .?AVbad_typeid@std@@    �X    .?AV__non_rtti_object@std@@          �            .   .   P�������������������T���������������X�uww   ���5      @   �  �   ����                     @�    @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                $~    ~   ~   ~   ~   ~!   �}   �}   �}   �}   �}   �}   �}   �}    �}   �}   �}   �}   �}   �}   �}   �}   �}   �}"   |}#   x}$   t}%   l}&   `}�&         �D        � 0        .                           �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
          �      ���������              �        ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (�         �� ��                     @� P� `� v� �� �� �� �� �� �� �� �� 
� � 0� D� `� ~� �� �� �� �� �� �� ��  � � ,� >� F� T� f� �� �� �� �� �� �� � &� 4� B� \� l� �� �� �� �� �� �� �� �� � � 4� D� R� `� v� �� �� �� �� �� �� �� 
� � 2� B� R� b� p� ~�                                                                                                     @� P� `� v� �� �� �� �� �� �� �� �� 
� � 0� D� `� ~� �� �� �� �� �� �� ��  � � ,� >� F� T� f� �� �� �� �� �� �� � &� 4� B� \� l� �� �� �� �� �� �� �� �� � � 4� D� R� `� v� �� �� �� �� �� �� �� 
� � 2� B� R� b� p� ~�                                                                                                     � DecodePointer � EncodePointer �GetCurrentThreadId  �GetCommandLineA �HeapAlloc GetLastError  �HeapFree  RtlUnwind IsProcessorFeaturePresent %WriteFile dGetStdHandle  GetModuleFileNameW  GetLocaleInfoW  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  �GetCurrentThread  EGetProcAddress  �Sleep ExitProcess oSetHandleCount  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �HeapSize  rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage 9LeaveCriticalSection   FatalAppExitA � EnterCriticalSection  -SetConsoleCtrlHandler ?LoadLibraryW  �HeapReAlloc bFreeLibrary �InterlockedExchange �RaiseException  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �GetUserDefaultLCID  GetLocaleInfoA  EnumSystemLocalesA  IsValidLocale �SetStdHandle  $WriteConsoleW � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �                 0  �              	  H   X  Z  �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel>
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPAD   D   �9d;u;�;�;�;<!<�<�<�<�=�=�=�=�=$>D>d>�>�>�>�>?4?T?q?�?�?      �   0$0Q0q0�0�0�01D1t1�1�1222G2�2�23A3a3�3�3�34$4D4t4�45'5=5\5�6888 8�8�8�8�9�9�9):D:}:�:�:�:;�;�;�;�;<<<N<g<�<�<=.=I=n=�=�=�=@>�>�>b?�?�?�?�?   0  H   0'0g01$1@1�1�1	2 2>2H2e2}2�2�2�2�23�3\4�4�4(7C7�7�9B:|:�:�;   @  L   Z1�1�1!2313�5�586t6�6�7]8�8�8�899+9I9f9|9�9�9�9�9�9:*;<<�>�>�> P  4   +0=0&2$525�5�586O6r6�6�7`8::�;�=6>|?�?�?�? `     w0�0�01141L12e2�34$4D4d4�4�4�4�455K5�5�5�56F6j6y6�6�6�6�6�6�677+7=7O7X7v7�7�7�7�7�788D8R8_8w8�8�8�8�8�8�89929H9d9v9�9�9�9�9�9::&:T:b:o:�:�:�:�:�:�:�:;&;B;X;t;�;�;�;�;�;�;<$<6<?<]<~<�<�<�<�<�<=='=9=K=]=o=x=�=�=�=�=�=>&>8>A>_>�>�>�>�>�>�>�>?4?P?b?t?}?�?�?�?�?�? p  �   040Q0q0�0�0�011+1G1`1q1z1�1�12262J2\2n2�2�23'383A3T3�3�3�344*4<4b44�4�4d5y5�5�5d6�6�6�6�6747Q7�7�798U8�8�899U9�9�9�9:8:T:t:�:�:;�;�;,<Q<�<�<�<=4=T=b=�=�=�=�=�=>1>D>d>�>�>�>�>�>�? �  �   ,0T041T1t1�1�1242d2�2�2�23D3�3�3-444;4B4I4P4W4^4h4r4y4�4�4�4�4�4�4�4�4�4�4�45%5]5n5546�6�8v9�9m:�:3;a;~;�;�;�<=5=u=�=>T>�>�>?�?�? �  �   010D0d0�0�0�0�0�0141d1�1�1�1�12!2D2t2�2D3t3�3�3�3414T4q4�4�4�4545d5�5�5�5.6r6�6�6�6�67D7q7�7�7�7�78D8t8�8�8�8949T9�9�9�9�9�9:A:P:t:�:4;a;t;�;�;�;<A<a<�<�<�<=!=A=d=�=�=�=$>T>�>�>�>?Z?�?�?�? �  �   010T0�0�0�0�0�01-1j1�1�12$2J2�2�23 3�34Q4e4z4�4�4�45S5v5�5�56$6D6�6�6@7�7�7�7�78I8s8�8�8�8�8939T9�9�9�9�9:4:T:�:�:�:;A;a;�;�;�;�;<d<�<�<�<=4==�=�=�=!>>>h>�>�>�>�>?,?L?f?�?�?�?�? �  �   0"0_0s0�0�0�01.1Q1k1�1�1�1{2�2�2�2,343Y3�3�5_8x8�8�89 9W9�9�9d;h;l;p;�;�;+<0<�<�<�<�<$=T=�=�=�=�=>D>�>�>�>�>?4?T?�?�?   �  �   0D0�0�0�0d1�1�1�1$2�23$3D3�3�3�3�34$4D4d4�4�4�4�4�4�45!545T5t5�5�5�5�5616T6q6�6�6�67$7D7d7�7�7�78!818D8d8�8�8�8�8�8!9?9d9�9�9�9�9%:=:L:q:�:�:�:�:�:	;;�;�;�;5<u<�<=5=u=�=�=5>�>�>%?e?�? �  p   0U0�0�0E1�1�152�2�23e3�34U4�4�4E5�5�556�6�6%7u7�78e8�8�859u9�9:e:�:;U;�;<U<�<�<E=�=5>�>�>%?u?�?   �  �   0e0�01U1�1�1U2�2�253�3�34�4�4!5q5�5!6q6�67q7�7�7�7�8�89!9A9a9�9�9�9�9�9:$:Q:t:�:�:�:�:;4;a;t;�;�;<!<A<a<�<�<�<=1=Q=t=�=�=>!>D>d>�>�>�>�>?$?D?d?�?�?�?�?�? �  �   040�0�0�0L1w1�1�1Q2�2�23�3�3�3A4^4v4�45#5�5�5�5!6D6�637\7�78,8T8�8�8$9�9�9�9K:�:�:A;g;�;�;A<g<�<,=�=�=�=n>�>�>?>?S?�?�?   �   0|0�0141Q1a1t1�1�1�12$2T2t2�2�2�2343Q3t3�3�34 4B4~4�4�4�455Q5q5�5�5�5�5�6�6�6�6�6�6747Q7d7�7�7�7�78D8t8�8�8�8�8�8949W9�9�9�9':b:�:�:�:N;\;�;�;�;�;<4<d<�<�<�<�<$=D=t=�=�=�=$>D>d>�>�>�>�>?$?6?Q?d?�?�?�?�?�?  �   0$0a0q0�0�0�01$1D1a1t1�1�1�1�1�1242T2t2�2�2�23$3A3T3t3�3�3�3�34d4�4�4�4�4545T5t5�5�5�5�56W6�6�67S7�7�78$8T8�8�8�8�89!919D9d9�9�9�9�9:-:f:�:�:�:�:;&;T;t;�;�;�;<<D<b<v<�<�<�<�<=4=T=�=�=�=�=�=>4>Z>�>�>�>�>�>�>?$?>?R?b?�?�?�?�?�?        0%0>0^0�0�0�0�011?1\1p1�1�1�1�1�12.2O2l2�2�2�2�2�23&3G3d3x3�3�3�34'4D4X4n4�4�4�4545T5t5�5�5�5�56$6A6T6�6�6�6�6747T7t7�7�7�7�78!848Q8d8�8�8�89$999K9T9e9{9�9�9�9�9�9:4:F:Y:l:�;�;�;[<�<�<�<�<�<=
====&=-=4=;=B=I=P=�>?$?D?a?t?�?�?�?�?   0 �   0$0T0t0�0�0�0141F1t1�1�1�12!2D2�2�243t3�3�3�3�3444T4t4�4�4�4545T5�5�5�5�5!6D6q6�6�6�67A7d7�7�7�7818Q8q8�8�8�8�8919Q9q9�9�9�9�9:1:;2;b;�;�;<E<�<�<=%=e=�=�=*>q>�>�>5?u?�?�?   @ �   0e0�0�0%1u1�1�12U2�2�2�2E3�3�34U4�4�4�4�45%5u5�5�526u6�67R7�7�7�78#8P8U8}8�8�8�89U9y9�9�95:Y:�:�:�:;?;x;�;�;<'<H<�<�<�<=V=�=�=>4>T>t>�>�>�>�>�>?%?3?T?e?s?�?�?�?�?   P (  0!010T0l0�0�0�0�0�0 11101T1l1�1�1�1�1�1�1
22+2=2a2q2�2�2�2�2343F3T3g3�3�3�34$4A4T4t4�4�4�45545T5t5�5�5�5�5�56$6D6d6�6�6�6�67$7D7^7u7�7�7�78#8>8U8m8�8�8�89%9=9T9�9�9�9�9 :(:<:�:�:�:;!;E;�;�;�;�;<$<D<d<�<�<�<�<=!=1=D=q=�=�=�=�=�=�=>#>1>@>a>�>�>�>�>�>??!?4?T?o?}?�?�?�?�?�? `   040T0t0�0�0�0�0'1@1Q1m1�1�1�1�1�1	242T2t2�2�2�2�233.3>3P3t3�3�3�3�3�3�34>4U4l4}4�4�4�4�4�45"565E5U5f5�5�5�5616D6t6�6�6�6�6�67$7D7d7�7�7�7�78$8D8d8�8�8�8�89$9D9d9�9�9�9�9 :D:d:�:�:�:�:;$;D;d;�;�;�;�;<$<D<d<�<�<�<�<=$=D=d=�=�=�=�=�=>1>D>a>q>�>�>�>�>�>
??D?d?�?�?�? p �   0"0�0�0�0T1t1�1�1�1�1�142Q2d2w2�2�2�23$3A3o3�3�3q4�4�4�4�4515D5t5�5�5�56$6D6t6�6�6�6747T7q7�7�7�7$898H8�8�8�89!9A9d9�9�9�9::A:�:�:;D;a;t;�=�=�=�=�>�>   � �   80q0�0�0�0111A1Q1a1�1�1�1�1$2D2g2u2�2�2�2�2313D3t3�3�4�455�5�6�6�6S7f7v7�7!8+8�9�9�9:4:T:t:�:�:�:�:$;D;d;�;�;�;�;<A<�<=   �    �8�8�9   � \   �3�34U4�4�4%5e5�5�56E6�6�6�657u7�7�7"8R8�8�8�8%9e9�9:E:�:�:;U;�;<e<�<�<5=?7?   � �   �1(2,20242823)3H3V3�3�34#4�4�4!5/5o5}5�6�6�6�6@7N7c7q7t8�8�8�8�899(9U9w9�9�9�9:2:�:�:�:�:�:�:�:;";3;F;Y;q;�;�;�;�;�;(<9<K<\<m<<�<�<�<�<$=1=7=c=j=�=�=�=�=�=>>> >$>(>1>T>�>�>$?V?   � T   0(0�0�0:4�4�4<6p6�677&7E7V7}7�78]8�9�:�:�:�:�:�:�:�:�:�:�:T;�<==m>v>�>�? � @   H1L1P1T1�1�1�1�1�1"2�2�2�2�2�5�5f6�;<�<!=/=�=�=�>>?o?�? � �   �0�041�1�1�1�1�1 222h2|2(3�3�3[4�4�435�5686<6@6D6H6L6P6T6X6\6`6d6v6�6�67�7�7�7�7�7?8W8p8�8�8�8�8�8�8&9>9S9g9�9�9�9�9�9:$:9:K:\:z:�:	;v;�;�<�<   � 4   &3�3n5�5�5�5O6b6�6�6�<�<�<�<F=X=l=�=�=�=�>     @   �2�2�2�2�2�23'3x3�3�344�5�5K6Z677�7�7�:�:�;�;<=%=  �   �1�12'2�2�2�3�3�4�4�7�7�7�7�7�7�7�7�7�7�7�7�7�7�788888%8p8�8,9D9K9S9X9\9`9�9�9�9�9�9�9�9�9�9�9�9::@:D:H:L:�:�:�:�:�:�:�:;7;i;p;t;x;|;�;�;�;�;�;�;�;�;�;J<==.=�=�=�=�=�=>>>>+>c>h>r>�>�>�>�>?<?B?H?]?�?�?�?   \   0C0�0�0�0.131<1K1n1s1x1�1�12202_2e2t2�2�2�203B3�3�3�34L5d5i5�7�7\8d8y8�8l;�;<   0 �   �1f24#4)45#506P6U6�6�6�6�7�7�78858�8A9;:d:v:�:�:�:�:;;2;:;@;N;�;�;�;�;�;><l<�<�<�=>?>Q>W>]>c>i>o>v>}>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????"?(?>?E?O?V?g?m?x?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @ \  0000(0J0_0�0�0�0�0�011/1U1�1�1�142<2�2�2�2�2�2�2�2�2�2�2�2�2�233 3(3.353;3B3H3P3W3\3d3m3y3~3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444?4E4]4�4�4�4�4�4�4�45 5,5e5n5z5�5�5�5�5�5�5�5 6�6�677-787=7O7Y7^7z7�7�7�7�7�7�7�7�7�728<8b8i8�8�8�8Y99�9�9�9�9:W:a:�:�:�:�:;(;V;y;;�;�;�;�;�;+<5<v<�<�<�<�<�<v>�>�>�>�>�>??.?V?�?�?�?�?�?�?   P x   00%0+01080A0^0�0�1�1�1�1N2�34(444<4D4P4y4�4�4�4�4�4	55�5�5�566%6+676=6Y7�7h8�8�9�:�:�:�:�:�:�:;;�;=�?   ` 8   0K0}0.1�1/2�3J5�9�9::#<=c=n=t=�=�=�=�>�>�>   p �   S0d0�0�0�0�0�0�0
11181B1U1y1�1�1�1h2�2�2=3�344.4@4[4c4k4�4�4�4�4�4�4�4�4
535D5X5�5�5;6�6R7�7�78#8\8�8�8�9�9�9�9�9�9�9�9�9::::@:�:�:;;�;�;<<�<�<	==�=�=	>>�>�>??�?�?   � �   0&02=2�2�3�4�4�4�4555595_5}5�5�5�5�5�5�5�5�5�5�5�5�5�5b6m6�6�6�6�6�6�6�67 7$7(7,7074787<7�7�7�7�7�7�8�8�8�:~<�<�<�<�<�<�<�<�<=#=)=7=J=]=�=�=>5>�>�>�>�>�>?$?U?�?�? � �   �0�0D1G2q2�2�3�3�3�3�3�3�3�3�3�3�3�3�3�344 424@4N4\4g4r4}4�4�4�4�4 5�6�6�6q7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�788(8	99 9&9/969=9F9N9T9Z9~9�9�97:�:0;E;�;<�<�<=9=J=�=>?n?�?   � �   1�1�1�1l2�2�2!303x3�34"4.4Y4h4�4�4�4 5�5�5�5
6r6�673787?7F7M7Z7c7�7�7�7�7�7�7�7�7�7�7"8H8N8Z8a8�8�8�8�8�8�8�8�8�89:9o9t9�9�9<:S:v:�:�:�:;;';x;�;�<�=
>>>o>z>�>�>�>�>	???"?,?G?[?q?�?�?�?   � �   000�0�01!1?1�1�1�12$2�233,3J3{3�3�34+4V4i4p4�4�4�4�4�4515T5q5�5�5�56#6\6v67*7N7�7�78-8=8�8�8�8�8�809=9F9f9a:�:�:;;9;D;^;�;�;�;�;<	<<<"<0<6<E<{<�<�<�<�<=-=9=S=\=�=�=�=�=�=�=)>;>`>|>�>�>�>�>?u?�?�?�?�?   � �   40U0j0�0�0�0�0�0�0)1.1D1i1�1�1�12;3 4)4E4[4�5�5Y6�6�6�6Y7�7838�8�8�9.:�:�:d;�;!<=,=�=�= >o>�>�>�>�>?'?8?O?X?�?�?�?�? � �   40d0�0�0�0u1�1�1�1�12_2�2�2�23-3M3l3�3�3	4V4m4�4	5{5�5�5�5l6�6d7�7�7>8}8�8&9�9�9�9�9�:�:F;c;{;�;�;"<�=�=�=�=>$>0>C>P>e>r>x>�>�>�>�>�?�?   � @  0I0Q0W0]0c0�0�0�0�0�0�0�0$1Q1g1�1�1�1�1�1�1�122I2`2v2�2�2�2�2�2333G3m3�3�3�3�34!4�4�4�4�4�4�4�4�4�4�45V5q5|5�5�5�5�56,6?6h6m6z6�6�6�6 77#707A7�7%818<9k9p9u9z9�9�9�9�9�9�9�9&:U:[:u:�:�:;N;�;�;�;�;�;�;�;�;�;�;<<<<%<3<8<@<F<T<Y<�<�<=;=@=G=L=S=X=f=�=�=�=^>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?	???'?b?|?�? � `   �1�1�1�1�2�2s3�344%4�4�4�4�4�4|5�5�5�5�5�5�56&636;6I677/7M7a7g7�;�;�<�=�=�=5>D>_>     l   t1j2�3A4m4�4r6�8�8�8�8�8�8�8�89�91:F:_:�: ;<;I;e;r;�;�;�;�;�;(<=<l<�<�<�<=<=r=�=	>\>�>�>E?_?h?�?�?  $   �0`1�1�1�2>�>-???Q?c?u?�?     �   �0�0�0�0�0"1�1�1�1�122'292K2]2o2�2�2�2J5�5�566$6*6;6C67#7C7I7�7�7�7�7�7�7(848u8�8G9":�:;);�;�;�;�;�;�;<j<�<>=;>�> 0 4   �01j1�1�12�2�2�2�2�4)5�5�5666)656@6<   @ H   V1�1�2�2�3g4�45�5�5�5V6m6�6*78&8�8�9P:V:�:�:;�;�;�;:=�?�?�?   P 8   �273�56W9[9_9c9g9k9o9s9w9{99�9�9\:;F;V;s;�;�; `    �37�9=<H?   p \   c2�5�5�5�5 6(6�67�7�7�8�8O9�:�;g<�<�<�<=�=�=>�>�>
??"?<?K?X?d?t?{?�?�?�?�?�?�?�? � d   0,0_0n0w0�0�0�02-2<2C2N2b3�3s6�78-8C8K8�8�9�9�9W:�:�:N;�;<v<4=F=X=�=�=�=�=�=>,>?>]>�>�? � \   =122#2-2X2`2�2�2�2�2�2�214L4]4}4�4�4�4:5v5�5<6_68J8�8�80999{9�9�9:\:e:~:�:�:;!; �    �0   � L   0"0&0*0.02060:0>0B0F0J0N0R0V0Z0^0b0f0j0n0r0v0z0~0�0�0�0�0�0�0�0(5   � d   r5v5z5~5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5&7>7�;�;�;�;�>�> ??�?�?�?�? � |   0"0:0Z0�0�0�0
171d1o1�1�1�1�12B2g2t2�2�2�23M3�3�3�3M4h4u4�4�4�5�56<6E6l6y6~6�6g7�7�7�78A8�8�8m9�9:8:T:p:�:a=�> � <   �1�1�1�1�12�2�2�233+4�4�45v5�5�5�8�9T;�;�;�;�=   � 0   3070;0?0C0G0K0O0Z2�23B3�34�4?;�=�=�=>   �   .2f2R5V5Z5^5b5f5j5n5�556?6W6�6�6�6t7z7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78
8888"8(8.848:8@8F8L8R8X8^8d8j8p8v8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 999999$9*9        �1�1 2C2u2�2�2�2     q3        �3�3�3�3�3�3 @ t   14444,7088><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? P l   004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�01 1014181<1@1D1H1�1�1�1�1�1�1h3l3�3�3�3�3�3�3�8�8�8 ` (  \1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12�2�2T4X4\4`4h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?   p D   �3�3�3�3�3�3�3�3�3�3�3�3`<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<   � �   0383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�6�6 �   |4�4�4�4�4�4�4�4�4�45550585<5@5H5`5x5|5�5�5�5�5�5�5�5�5�5�5�5666(686<6L6P6X6p6�6�6�6�6�6�6�6�6�6�6�6�6�6777,70747<7T7d7h7x7|7�7�7�7�7�7�7�7�7�7�7�788808@8D8T8X8\8d8|8�8�8�8�8�8�8�8�8�8�8�899 9094989@9X9\9t9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :8:H:L:\:`:d:h:p:�: � �   �1222 2(20282@2H2P2\2�2�2�2�2�2�2�2�2�2�2�2�2�23$303P3\3|3�3�3�3�3�34(4H4h4�4�4�4�4�4�4585@5D5\5`5|5�5�5�5�5�5�5�5�56 6(6X6`6d6|6�6�6�6�6�6�6�6�6�6�6�677,707P7p7�7�7�7�7808P8l8p8�8�8�8�8�8�8�8989X9t9x9�9�9�9�9 : :@:L:h:�:�:�:�:   � @   0080`0�0�0�0�0 1$1H1d1�1�1�1222222 2$2(2,2�34X8X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;(;8;H;X;|;�;�;�;�;�;�;�;�<�<�<�<=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�= � D   t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      