MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       #�p\B�#\B�#\B�#`�#]B�#�^�#FB�#`�#6B�#\B�#B�#>]�#_B�#`�#qB�#�b�#]B�#Rich\B�#                        PE  L �LH        � !    �      xv                               �                              �/ G   �* (                            � �                                                     �                           .text   �                         `.rdata  �                       @  @.data   �d   0  P   0             @  �.reloc  �"   �  0   �             @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���   �lySU��$�   V�ًHHW�T$lUR�\$<�QH�   ��ly��$�   �HHj h'  U�Qx�����l$8u_^][���   � �SR�4 ���D$$��u_^][���   � �C3���v!�ly��$�   VU�HDVR�QD�C��F;�rߋC�{@���D$,    �8  ��|  �|$����  ��$�   j QP��$  ��$�   RP�5 ���D$0��t=�K3���v%��D$0�lyVP�D$,�QDVP�RD�C��F;�rݍL$0Q��5 ���(�C3���v�ly�L$$VU�BDVQ�PD�C��F;�r�7��$�   �D$  �?�D$  �?�H/ �ly��$�   QV�B@�P`����$�   ��$�   R�\/ ��$�   �/ j h�  ��$�   �0 ���\$j h�  ��$�   �t0 ���\$ j h�  ��$�   �[0 �\$(j h�  ��$�   �D0 �D$(�� ����@u�� �t$(�\$�� ����@u�� ���\$�G�3�����m  ��|$�G��L$4�ly�D$t    ���q4�D$p    �D$l    ��Ǆ$�       ����D$|    �D$x    Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       �BD�S�L$lQ�L$(RQ�P<�D$x�L$�   �t$x�|$H�ly�D$$��\$H�D$T�L$�D$$�L$HQ��$  �\$X�D$d�L$ �D$(�\$d�D$p�L$ �D$(�\$p�D$P�L$$�D$0�\$P�D$\�L$$�D$0�\$\�D$h�L$$�D$0�\$h�D$t�L$$�D$0�\$t�BD�SRQ�P@�T$4��E;j�������\$4����$�   �t- �l$8�D$,�K�ǀ  @;��|$�D$,������D$$P�(3 ���   _^][���   � ���SVW���&: �~���; ��> �^,�G��� !�t; ��> �C� !hL0���� ��% h@0����% �D$_�F@��^[� ���������SV��W�~,�_S�> �����    �O; �~�_S�s> �����    �3; ���9 �D$t	V�_? ����_^[� ����V��W�~W�3> �����    ��: �D$t	V�&? ����_^� ��������������V����8 ��t_j j j ���d8 ��tN�D$j�NPQ���D$   �D$    ��7 �T$j�F,RP���D$   �D$    �7 �   ^���3�^��Ð������������V���e8 ��u^��ËF@SUW3��D$   W�|$���  jh�� j�T$ QR���6 �F@�D$   �|$W���  �T$QR���5 �F@9�$  u2W�D$�   WP�Ή\$�|$ �5 �L$WQ�Ή\$�|$�=5 � �D$   �|$��   W�D$RP���[5 �N@�   �\$�|$���  W�D$RP���75 �F@9�   tfW�L$jQ���D$   �|$ �5 W�T$WR���D$   �|$ ��4 W�D$WP���D$   �|$ ��4 W�D$   �|$W�L$�<  9�  tgW�T$WR���D$   �|$ �4 W�D$jP���D$   �|$ �4 W�L$WQ���D$   �|$ �o4 W�T$W�D$   �|$R��   9�  tdW�D$WP���D$   �|$ �54 W�L$WQ���D$   �|$ �4 W�T$jR���D$   �|$ � 4 W�D$W�D$   �|$P�bW�L$WQ���D$   �|$ ��3 W�T$WR���D$   �|$ �3 W�D$WP���D$   �|$ �3 W�D$   �|$j�L$Q���3 �V@9��  tFW�D$jP���D$   �|$ �\3 �L$jQ�Ή\$�|$�3 �T$j�D$   �|$R�'�D$WP�Ή\$�|$��2 �L$W�D$   �|$Q����2 �V@9�  tLW�D$jP���D$   �|$ ��2 �L$j�   Q�Ήl$�|$�2 �   �T$j�\$�|$R�-�D$�   WP�Ήl$�|$�R2 �   �L$W�\$�|$Q���82 �V@9�  t(W�D$jP�Ήl$�|$ �V2 W�L$W�\$�|$Q�&W�T$WR�Ήl$�|$ �/2 W�D$j�\$�|$P���2 �N@�D$   �|$W��  �D$RP����1 �N@�D$   �|$W��  �D$RP����1 �N@9��  t0W�T$jR���D$   �|$ �1 �D$j�D$   �|$P��L$W�D$   �|$Q���>1 �V@�D$   �|$W���  �L$PQ���[1 �V@�	   �l$�|$���  W�L$PQ���71 �V@�
   �\$�|$���  W�L$PQ���1 �V@9��  tBW�D$jP���D$   �|$ ��0 �L$jQ�Ήl$�|$�0 �T$j�\$�|$R�#�D$WP�Ήl$�|$�q0 �L$W�\$�|$Q���\0 �V@�D$   �|$W���  �L$PQ���y0 _][�   ^��Ð������������D$���  HS�   V;�W����	  3Ɋ��% �$�d% �T$��$�  3�RP��Ǆ$�     ��$�  ��0 ����	  9|$tN��$�   jQ��Ǆ$     ��$  �/ �T$,jR���D$4   �|$8�/ _^�   [���  � ��$l  WP��Ǆ$t     ��$x  �N/ �L$<WQ���D$D   �|$H�5/ _^�   [���  � �T$��$  3�RP��Ǆ$     ��$  �,0 ����  9|$tN�L$LjQ���D$T	   �|$X��. ��$�  jR��Ǆ$�  
   ��$�  �. _^�   [���  � �D$\WP���D$d	   �|$h�. ��$  WQ��Ǆ$$  
   ��$(  �e. _^�   [���  � �T$�D$l3�RP���D$t   �|$x�e/ ����  9|$t4��$|  jQ��Ǆ$�     ��$�  �. _^�   [���  � �T$|WR��Ǆ$�      ��$�   ��- _^�   [���  � �D$��$,  P3�Q��Ǆ$4     ��$8  ��. ���S  9|$�I  W��$�   WR��Ǆ$�      ��$�   �- W��$�  WP��Ǆ$�     ��$�  �- W��$�   WQ��Ǆ$�      ��$�   �`- _^�   [���  � �T$��$<  3�RP��Ǆ$D     ��$H  �. ����  9|$��  W��$�   WQ��Ǆ$�      ��$�   ��, W��$�  WR��Ǆ$�     ��$�  ��, W��$�   WP��Ǆ$�      ��$�   �, _^�   [���  � �L$��$L  3�QR��Ǆ$T     ��$X  �c- ����  9|$��  W��$�   WP��Ǆ$�      ��$�   �>, W��$�  WQ��Ǆ$�     ��$�  �, W��$�   WR��Ǆ$�      ��$�   ��+ _^�   [���  � �D$��$\  P3�Q��Ǆ$d     ��$h  �, ���7  9|$�-  W��$�   WR��Ǆ$�      ��$�   �+ W�D$WP���D$    �|$$�p+ W�L$ WQ���D$(   �|$,�V+ _^�   [���  � �T$�D$$3�RP���D$,   �|$0�, ����  9|$tA�L$4jQ�Ή\$<�|$@��* �T$DjR���D$L   �|$P�* _^�   [���  � �D$TWP�Ή\$\�|$`�* �L$dWQ���D$l   �|$p�i* _^�   [���  � �T$�D$t3�RP�Ή\$|��$�   �j+ ����  9|$��  W��$�   WQ��Ǆ$�      ��$�   �E* _^�   [���  � �T$��$�   3�RP��Ǆ$�      ��$�   ��* ����  9|$�z  W��$�   WQ�Ή�$�   ��$�   ��) _^�   [���  � �T$��$�   3�RP��Ǆ$�      ��$�   ��* ��t"�N@�T$���  �F@9��  u
ǀ�     �F@��$�      Ǆ$�      PQ�Ή�$�   �B* �V@��$�   ���  ��RPǄ$�      ��$�   �* �N@��$�   ���  Ǆ$�      QR�Ή�$�   ��) �F@��$�   �  Ǆ$�      PQ�Ή�$   ��) �V@��$  ���  ��RPǄ$     ��$  �) �N@��$  ���  Ǆ$     QR�Ή�$   �l) �F@��$$  �  Ǆ$$     PQ�Ή�$0  �B) �V@��$4  ���  ��RPǄ$<  	   ��$@  �) �N@��$D  ���  Ǆ$D  
   QR�Ή�$P  ��( �F@��$T  �  Ǆ$T     PQ�Ή�$`  ��( �V@��$d  ��   ��RPǄ$l     ��$p  �( �N@��$t  ��  Ǆ$t     QR�Ή�$�  �l( �F@��$�    Ǆ$�     PQ�Ή�$�  �B( �V@��$�  ��  ��RPǄ$�     ��$�  �( �N@��$�  ��  Ǆ$�     QR�Ή�$�  ��' �F@��$�    ��$�  PQ�Ή�$�  ��' �V@��$�  ��  ��RPǄ$�     ��$�  �' �N@��$�  ��  Ǆ$�     QR�Ή�$�  �p' _^�   [���  � �I " � l < � � � 5 �  8! �! P%  	
��������D�L$ SV�t$PWV�\����G ��3�SS�Gj����  �O8���  �W<���  �GD���  �OH���  �WL���  �G@���  �OP���  �WT���  �GX���  �O\��   �W`��  �Gd��  �Oh��  �Wl��  �Gp��  �Ot��  �Wx��  ���   ���  ���   ��   j��L$�
( ��uF�T$HR�, ���L$8�\$H�L) �D$4P�r, ���L$$�\$4�2) �L$�' _^3�[��DË��  �O���  �W8���  �G<���  �OD���  �WH���  �GL���  �O@���  �WP���  �GT���  �OX��   �W\��  �G`��  �Od��  �Wh��  �Gl��  �Op��  �Wt��  �Gx���  ���   ��$  ;�t��   ���   �� ���  ;Ë��  tB;Ë��  t;�tǆ�     �hǆ�     �\;�tǆ�     �Lǆ�     �@;Ë��  t;�tǆ�     �&ǆ�     �;�tǆ�     �
ǆ�     �D$HP��* ���L$8�\$H�' �L$4Q��* ���L$$�\$4�' �L$�& _^�   [��DÐ�������������$�lySUVW�|$8�L$h�  �HHW���   ���ϋ��� �؅���   �+ �L$�D$8�%- �L$8j W��+ ��uFh�0�L$(�. �T$$R�0 ���L$$��. �L$��, �D$8P�~+ ��3�_^][��$� 3���~%�L$j �.Q�L$@RW�t, ��t1�|$ PF;�|ۍL$�, �T$8R�1+ ��_^]�   [��$� h�0�L$(�. �D$$P�'0 ���L$$�+. �?�T$h\0�L$(ǂ$      ��- �D$$P�3) ���L$$������- ���v����L$�!, �L$8Q�* ��3�_^][��$� ����������@SU�L$VW�L$� �\$T���9  �ly3�Wh�� �HHS�|$`�Qx������tu�L$(�v �ly�L$(QV�B@�P`���T$(�L$<R� �L$(�� �D$<�L$P�� �L$<� Wh�  �L$�4 ����tj h�  �L$� �D$T���� �ly�苑�   ���R=�  u/��u+��t��u"�D$X��t�t$S��������tu��$  ��tS�t$X��u�   ���u3��D$T��u�ly�ˋ��   �R4�L$VP������ly�ˋ��   �R(�؅�������L$�� _^]�   [��@� �L$�� _^]3�[��@� ����������VW�|$����  SU�ly�ϋ��   �R=�  ��   �lyj h�  W�HH�Q|�ly��h�  W�BH���   �lyh�  W�؋QH���   ���   ���  ��Ѕɉ��   ��tÉ��   ���  ��u
���  ��tD��~@���  �E��t���   ��t���   �(;ht��t���   ��t���   ��Kuɡly�ϋ��   �R4P��������ly�ϋ��   �R(���������][_^� ��������������xSUVW�L$t�� �L$d�g* ��$�   3ۋ�$�   ���L?��\  ��\  �D$�n\���\  �D$��\  �D$;���  �?�D$D  �?�D$H  �?�D$L  �?�] ��\  ��\  �F@  �B�FD  �B�FH��N�N�^�^�^�^�F�F �F$�F(�F,�^0�^4�^8�F<�^P�^L�^T�^X�I  �ly�ϋ��   �R=G  �.  �lySW�HT�Q0�����  �lySW�BT�P,���L$PQ���W/ P�L$x�] �L$P�D �D$4  �?�T$4�D$8  �?�D$8�T$D�D$<  �?�L$<�T$D�D$HR�D$T�L$Ph�  P��$�   �I �h  �?�L$8h�  �P�L$|�T$@�@�D$D�� �D$4�ɍL$$��D$8���^�D$<���^���( P�L$Th�  Q��$�   �V P�L$h�<) �L$P�) �L$$��( jh�   U�L$p�9* �   �nP��   �lyjW�BT�P0������   �L$�', �lyjW�QT�R,���L$PQ���. P�L$x� �L$P� Sh�  �L$|� �^�T$S�D$TRP�L$0�D$\�  �\$`�\$d��, P���- �L$$��, �L$�V, �^H�L$�, �lyUW�QT�R0�����  �lyUW�HT�Q,���T$P��R�u- P�L$x�{ �L$P�b �D$$    �D$$�D$(    �L$(�D$D�D$D�L$HP�L$T�D$0    �T$0h�  Q��$�   �T$X�g �h  �?�T$8h�  �H�L$@�L$|�P�T$D�  �D$4�ɍL$$�^�D$8���^�D$<���^����& P�D$Th�  P��$�   �s P�L$h�Y' �L$P� ' �L$$�' j��\  h�   P�L$p�P( �nL�lyjW�QT�R0�����2  �nT�lyj	W�HT�Q0�����  �lyj	W�BT�P,���L$PQ���), P�L$x�/ �L$P� �D$$    �T$$�D$(    �D$(�T$D�D$,    �L$,�T$D�D$HR�D$T�L$Ph�  P��$�   � �h  �?�L$8h�  �P�L$|�T$@�@�D$D� �D$4�ɍL$4�^ �D$8���^$�D$<���^(���~% P�L$Th�  Q��$�   �' P�L$h�& �L$P��% �L$4��% j��\  h�   P�L$p�' �nX�lyjW�BT�P0������   �lyjW�QT�R,���L$PQ����* P�L$x�� �L$P�� �L$4��$ P�T$Th�  R��$�   � P�L$h�l% �L$P�3% �L$4�*% �D$jh�   P�L$p�e& �lyjW�QT�R0������   �lyjW�HT�Q,���T$P��R�^* P�L$x�d �L$P�K �L$4�B$ P�D$Th�  P��$�   �� P�L$h��$ �L$P�$ �L$4�$ �L$jh�   Q�L$p��% �lyjW�BT�P0������   �lyjW�QT�R,���L$PQ����) P�L$x�� �L$P� �L$4�# P�T$Th�  R��$�   �O P�L$h�5$ �L$P��# �L$4��# �D$jh�   P�L$p�.% �L$d��# �L$t�L _^][��xÐ�����P  SUV��W��$�   � ��$�   � �ly�V3�HU��UR��$�   ��$�   �l$P��H  ��;ŉD$��  �NU��QP�4 �ly�NUU�B��Q��H  ��;ŉD$u2h<2�L$d��" P�= ���L$`�# �T$R� ���1  �NU��QP�� �N�n�lyU���BUQ��H  ��;ŉD$u<h(2�L$d�" P�� ���L$`�" �T$R�Q �D$ P�G ����  �NU��QP�a �ly�NUU�B��Q��H  ��;ŉD$$uFh2�L$d� " P�j ���L$`�>" �T$R�� �D$P�� �L$$Q�� ���J  �VU��RP�� �ly�VUU�H��R��H  ��;ŉD$uPh�1�L$d�! P�� ���L$`��! �D$P�n �L$Q�d �T$$R�Z �D$0P�P ����  �NU��QP�j �ly�NUU�B��Q��H  ��;ŉD$(uZh�1�L$d�)! P�s ���L$`�G! �T$R�� �D$P�� �L$ Q�� �T$(R�� �D$4P�� ���?  �NU��QP�� �ly��$p  Uh�� �BHS�Px����;�t}��$�   ��	 �ly��$�   PW�Q@�R`����$�   Q��$�   ��	 ��$�   �
 ��$�   ��$�   R�
 ��$�   ��	 Uh�  ��$�   �
 ��$�   �lyUh�� S�HH�Qx����;�tz��$�   �8	 �ly��$�   QW�B@�P`����$�   ��$�   R�L	 ��$�   �	 ��$�   ��$�   P�|	 ��$�   �`	 Uh�  ��$�   �
 �D$x3��ly��PG�QHh)  S��$�   �Rx�������  �ly�͋��   �RxP��$�   �! ��$�   �� ��u��$�   �e �3ۉ\$ �ly��P��$h  �QHh�  PC�Rx��������   j ���� ��$�   �D$H� �ly��$�   PW�Q@�R`����$�   Q��$�   �. ��$�   �b ��$  �V P��$�   h�  R��$�   ��	 ��$�   �0 ��$  � ��$�   � ��t��$�   ��$�   P�p ��u��$�   �p ������$�   �D$    �W ��$�   3���~u��$�   � ���  P��$   QR��$�   �b	 ��$�   � ��$  ��$�   P�� ��u��$  �� G;�|���D$ ��$  �D$ �� �\$x3���~c�L$L�B ���  P�T$dQR��$�   �� �L$L� �D$`��$�   P� ��u�L$`� G;�|���D$ �L$`�D$ �h ���
 �   �T$4�L$@�L$<�L$0�L$8�L$,�D$\QRj ���u# ���G  �\$ �|$4�D$,;��  �Ë�����D$p�Ã��D$t��t\�D$�<� uR�D$H��tJ�ly���   ���R=G  u2�D$0��t�F�D$0    @�F�D$��   �N�T$����A��D$p3�;�t<�D$9�u39L$@t���  �L$@�� ���  �VB�V��   �F�T$$��� 9L$tt<�D$9�u39L$<t���  �L$<��@���  �VB�V��   �F�L$(��� �D$,G;������L$8�T$,��A�L$8�L$4RQ�L$dP�." ���������$�   �� ��$d  �|$|�����F3Ʌ�v8�T$�<� u�D$� �D$�<� u�D$$� �T$�<� u�D$(� �FA;�rȋVj Bj �V�ly�Q�@����P��H  ���F@��u h�1�L$P� P�e ���L$L�'  �N3�U�I����QP� �F��3�;�vY3��T$��;�t4�lyU���QUP��H  �N@����9x  �V@9�:x  ��   �
�F@��8x  �FC�ǀ  ;�r����  �nQ�L$P�{ P�F�N@�@������`  � �L$L� 9��  t�V@���  RP�n������VUBU�V�ly�Q��    +���Q��H  ��;ŉF8u|h�1�L$P�� P�F ���L$L� �T$R�� �D$P� �L$ Q� �T$(R� �D$4P� �L$<Q�  h�1�L$P� P�� ���L$L�  �NU��    +���RP� �F��3�;�vM3��D$$��;�t.�lyU���QUP��H  �N8���D9�V89l:�l  ��F8�l8�FC��;�r���$h  �����3����It�   �|� u�D$D@�x�;�r�L$D3�h�1�^�,��$  �� PU��$  �� �T$PPR�{ ���V8P�F��    +ȍ��  �L$L�� ��$�   � ��$  � �FS@S�F�ly�Q��    +���Q��H  ��;ÉF<��   h�1�L$P�> P� ���L$L�\ �T$R� �D$P�� �L$ Q�� �T$(R�� �D$4P�� �L$<Q�� ����$�   � ��$�   � _^]3�[��P  � hl1�L$P� P� ���L$L��  �NS��    +���RP� �F��;�vW3��D$(����t2�lyj ���Qj P��H  �N<���D�V<�D���K  ��F<�D    �FC��;�r�3�hd1��$  �^� PU��$  � �L$PPQ�� ��P�F��    +ЋF<���F �L$L� ��$�   � ��$  �� �N�T$��SQR�� �F�L$ ��SPQ� �V�D$0��SRP� ��$��$<  �0 ��$,  �$ 3��\$D�ly��P��$h  �QHGh)  P��$�   �Rx���;��7  �ly���   ���RxP��$�   �� ��$�   �� ����   ��$�   �/ �hD1�L$P�� P�9 ���L$L� �L$Q� �T$R� �D$ P� �L$(Q� �T$4R� �D$<P� ����$�   �B�  ��$�   �6�  _^]3�[��P  � ��$d  3��|$ �ly��Ph�  �QHSG�Rx���D$,���,  j ��� ���D$Ht�ly�L$H���   �R=G  t0�D$D��u(h1�L$P� P� ���L$L�# �D$D   ��$�   ��  �ly��$�   R�H@�D$0P�Q`����$�   Q��$P  � �  ��$�   �T�  ��$�   �H P��$�   h�  R��$X  ���  ��$L  �"�  ��$�   � ��$�   �
 ��t��$�   ��$�   P�b ��u��$�   �b �������$�   �D$    �I ��$�   3���~p�L$`� ���  P��$  QR��$�   �W�  P��$@  �: ��$  �� �L$`�� ��$<  ��$�   P�� ��uG;�|��
�D$ �D$ �\$x3���~v��$�   �6 ���  P��$   QR��$�   ���  P��$0  � ��$  � ��$�   �u ��$,  ��$�   P�Q ��uG;�|��
�D$ �D$ �����  �   �T$\�L$8�L$<�L$4�L$@�L$0��$�   QRj ���V ����  �|$\�D$0;���  �D$ ���ȋЃ�������$�   �T$p�D$t�����$�   ���  �D$�<� �  �l$H����   �ly���   ���R=G  ��   �D$4��t���  �F�ɀ@���  �F�ly�͋��   �RxP�F�@���F@����`  �w �F�@���F@�L$,����|  �F�N@�@�����PU�������D$4    �N4�V�T�F�@���F@���p  ��x  �<��F�@���F@����p  ��p  A��L$��   �D$p����   �T$�<� ��   �D$8��t-�n��$<  EQ�ŉn��    +ЋF8��� �D$8    �N4�V�T�F�V8��    +ȍ��L��P�<��F�V8��    +ȍD��L�A��D$��   �D$t����   �L$�<� u~�D$<��t+�F��$,  @R�V<�F��    +ȍ��
 �D$<    �F4�N�L�F��    +ЋF<�L����P�<��F�V<��    +ȍD��L�A��D$��   �D$0G��P;�������L$@�T$\��A�L$@�L$0Q��$�   RP� ���?�����$�   �A �|$|3������~�V�N�FGBA�~�N3�;ÉV��   3�3��V$׋j;j�V4t
�DL   ��DL   �V4��V4�\�V4�L�T$9�u"�V4�\�V@��p  ��x  ���V@��p  �T$9�u�V4�\�V8�j�R���V8�B�T$9�u�V4�\�V<�j�R���V<�B�VA����P;��I���9��  �A  3�ly��P��$h  �QHh�  PE�Rx�؃����  j �����  ����tǋly���   ���R=G  u���$�   ���  �ly��$�   RS�H@�Q`����$�   ��$L  P��  ��$�   �7�  ��$�   �+ P�L$dh�  Q��$X  ���  ��$L  ��  ��$�   �| �L$`�� ��uU���  �πʀ���  �ly���   �Px�N@P��`  �p �N@��|  �V@RW���  ǆ�     �������L$`� ��������  ��u�F@Pj ��������L$Q�	 �T$R�	 �D$ P�	 �L$(Q�|	 �T$4R�r	 �D$<P�h	 ����$,  � ��$<  � ��$�   ��  ��$�   ��  _^]�   [��P  � �����$SUVW�|$8��3�ωnL��  ;ŉF u_^]3�[��$� �����  ��;�u0h\2�L$(�� �D$$P� ���L$$� _^]3�[��$� �ly�F UU�Q��P��H  ��;ŉFLuhP2��  ��_^]3�[��$� �N U��QP� �F �~L��;ŉl$�Z  �\$��\$���� �S��lyj ��   j �HS�l$,�T$(��H  ���G��t��lyj j S�B��H  ���G���m����lyj j S�Q��H  3Ƀ�;��G�I����D$3�;���L$8�L$��  �D$� ������   @�d  ������X  �   ����I  ����n4#Ë؋��%�������͋)��   �)�l$�i���   @�  ������  �$��N �L$8��u=�^$�o������\� �^H��t
�o��\� �^0��t
�o��L� �D$8   B�N$�_���L���NH��t
�_�L���N0����  �_�D�q  �L$8��u@�^$�o�����\�\� �^H��t�o�\�\� �^0��t�o�L�L� �D$8   B�N$�_���L���NH��t
�_�L���N0���   �_�D��   �L$8��u@�^$�o�����\�\� �^H��t�o�\�\� �^0��t�o�L�L� �D$8   B�N$�_���L���NH��t
�_�L���N0����   �_�D�t�L$8��u@�^$�o�����\�\� �^H��t�o�\�\� �^0��t�o�L�L� �D$8   B�N$�_������NH��t	�_����N0��t	�_���B�l$ ;�}�L$�D$A;ȉL$�o����l$ �D$�T$�o�N �� @��;��D$�T$�����_^]�   [��$� IL �L FM �M SVW����  �~��� �g �^,�G��� !��  �O �C� !hL0���H!�d�  h@0���X�  �D$_�F@��^[� ���������3�Ð��������������V�����  ��t_j j j/���t�  ��tN�D$j�NPQ���D$   �D$    ���  �T$j�F,RP���D$   �D$    ���  �   ^���3�^��Ð������������V���u�  ��u^��ËF@W3��D$   W�|$��4  jh�� j�T$QR����  �F@�D$3   �|$W��L  �T$QR�����  �F@�D$4   �|$W��P  �T$QR����  �F@�D$5   �|$W��T  �T$QR����  �F@�D$6   �|$W��X  �T$QR���a�  �F@�D$7   �|$W��t  �T$QR���>�  �F@�D$8   �|$W��x  �T$QR����  �F@�D$9   �|$W��\  Q�T$��R���  �F@�D$2   �|$W��`  �T$QR�����  �F@�D$1   �|$W��d  �T$QR����  �F@9�8  t0W�L$jQ���D$@   �|$��  W�T$W�D$A   �|$R�.W�D$WP���D$@   �|$�]�  W�L$j�D$A   �|$Q���B�  �F@9�@  ttW�T$jR���D$<   �|$��  W�D$WP���D$=   �|$��  W�L$WQ���D$>   �|$���  W�T$WR���D$;   �|$���  _�   ^���9�D  ttW�D$WP���D$<   �|$��  W�L$jQ���D$=   �|$��  W�T$WR���D$>   �|$�l�  W�D$WP���D$;   �|$�R�  _�   ^���9�H  ttW�L$WQ���D$<   �|$�%�  W�T$WR���D$=   �|$��  W�D$jP���D$>   �|$���  W�L$WQ���D$;   �|$���  _�   ^���W�T$WR���D$<   �|$��  W�D$WP���D$=   �|$��  W�L$WQ���D$>   �|$�}�  W�T$jR���D$;   �|$�b�  _�   ^��Ð�������D$��  HV��@W����  3Ɋ�lY �$�LY �T$��$�   3�RP��Ǆ$�   @   ��$�   ���  ���b  9|$�X  W�L$$WQ���D$,A   �|$0���  _�   ^��  � �T$��$�   3�RP��Ǆ$�   A   ��$�   ��  ����  9|$��  W�L$4WQ���D$<@   �|$@�q�  _�   ^��  � �T$��$�   3�RP��Ǆ$�   <   ��$�   �)�  ����  9|$��  W�L$DWQ���D$L=   �|$P��  W��$�   WR��Ǆ$�   >   ��$�   ���  W�D$TWP���D$\;   �|$`���  _�   ^��  � �L$��$   3�QR��Ǆ$  =   ��$  ��  ����  9|$��  W�D$dWP���D$l<   �|$p�l�  W��$�   WQ��Ǆ$�   >   ��$�   �I�  W�T$tWR���D$|;   ��$�   �,�  _�   ^��  � �D$��$�   P3�Q��Ǆ$�   >   ��$�   ���  ���U  9|$�K  W��$�   WR��Ǆ$�   <   ��$�   ��  W��$�   WP��Ǆ$�   =   ��$�   ��  W�L$WQ���D$;   �|$ ��  _�   ^��  � �T$��$  3�RP��Ǆ$  ;   ��$  �:�  ����  9|$��  W�L$WQ���D$$<   �|$(��  W�T$,WR���D$4=   �|$8��  W�D$<WP���D$D>   �|$H���  _�   ^��  � �L$�T$H3�QR���D$P   �|$T���  ��t�F@�L$��4  �V@�D$X��d  ��RP�D$`1   �|$d�x�  �N@�T$h��`  �D$h2   QR�Ή|$t�V�  �F@�L$xL  �D$x3   PQ�Ή�$�   �2�  �V@��$�   ��P  ��RPǄ$�   4   ��$�   ��  �N@��$�   ��T  Ǆ$�   5   QR�Ή�$�   ���  �F@��$�   X  Ǆ$�   6   PQ�Ή�$�   ��  �V@��$�   ��t  ��RPǄ$�   7   ��$�   ��  �N@��$�   ��x  Ǆ$�   8   QR�Ή�$�   �\�  �F@��$�   \  Ǆ$�   9   PQ�Ή�$�   �2�  �V@��$�   ��8  ��RPǄ$�   @   ��$�   ��  �N@��$�   ��@  Ǆ$�   <   QR�Ή�$  ���  �F@��$  D  Ǆ$  =   PQ�Ή�$  ��  �V@��$  ��H  ��RPǄ$   >   ��$$  ��  _�   ^��  � �I �V ^V oT U �U �S T 9Y  �����D�L$ SV�t$PWV������G�  ��3�SS�Gj���4  �O��8  �W��@  �G��D  �O ��H  �W$��L  �G(��P  �O,��T  �W0��X  �G4��\  �O8��t  �W<��x  �GD��h  �OH��p  �WL��|  �G@���  �OP���  �WT���  �GX���  �O\���  �W`���  �Gd���  �Oh���  �Wl���  �Gp���  �Ot���  �Wx���  �G|��`  ���   ��d  j��L$��  ��uF�T$HR�>�  ���L$8�\$H���  �D$4P�$�  ���L$$�\$4���  �L$�k�  _^3�[��DË�4  �O��8  �W��@  �G��D  �O��H  �W ��L  �G$��P  �O(��T  �W,��X  �G0��\  �O4��t  �W8��x  �G<��h  �OD��p  �WH��|  �GL���  �O@���  �WP���  �GT���  �OX���  �W\���  �G`���  �Od���  �Wh���  �Gl���  �Op���  �Wt���  �Gx��`  �O|��d  ���   �e�  �D$HP���  ���L$8�\$H��  �L$4Q���  ���L$$�\$4��  �L$��  _^�   [��DÐ�������������H  SUV��W�L$��  �L$<�� �NP�J�  h�3�L$$���  ���  P��� �L$ ���  �D$ ��P�y P�L$��  �L$ ���  j�L$\h   Q�L$��  �T$XR�G�  �����L$ W�x�  P�L$���  �L$ ��  �D$�L$ P�G P�L$@� �L$ � �L$<Q���h ���nt��S�J ���c�  ����  ���  Wh�3S�y ���NdS�-�  �H3���3�S���+��ы������ʃ�����  �,3���3�S���+����������ȃ������  ��2���3�S���+��ы������ʃ�����  ��2���3�S���+����������ȃ�����  ��2���3����+�S�ы������ʃ����[�  ��2���3�S���+����������ȃ����1�  ��2���3�S���+��ы������ʃ�����  ��2���3�S���+����������ȃ������  �H3���3�S���+��ы������ʃ�����  ���L�  �L$<���  �L$��  _^][��H  Ð��������������U������   SUV��WhT4�L$$�\$�,�  P��  ���L$ �J�  �C�k@���D$    ��  j�D$4h   P��`  �m�  �L$0Q��  ���KP�D$P��  ����  �P4����Ü  ���+��D$�ы���S���ʃ��pt�����  �L$QhD4S�� ����S��  �ET��t(�E@�x!���MD�$h<4S�� ����S�|�  �E�� ����@uD�E�-p!���$h44S� ����S�G�  �EH���$h,4S�s ����S�(�  � 4���3�S���+��D$�ы������ʃ��pt�����  �EL��t1�E���$�E���$�E���$h4S�
 �� ��S��  �E���$�E���$�E ���$h 4S�� �� ��S��  �EX��t1�E(���$�E$���$�E ���$h�3S� �� ��S�V�  ��\  ��\  ��tPh�3S�z ����S�/�  �M\�E\��tPh�3S�Y ����S��  ��\  ��\  ��tPh�3S�2 ����S���  ��\  ��\  ��tPh�3S� ����S���  ��\  ��\  ��tPh�3S�� ����S��  ��\  ��\  ��tPh�3S� �L$ ����tS�m�  �\$�Kt��  �D$�K�ŀ  @;��D$����_^][��]Ð����������������  SUVW�����̍�  ���   P���  ����  3�;��   h   h�p�Ή_���  ��tZ��p<#t<<nu8�L$(Qhl4h�p�U ����uh�p�A�  �����   P��  �Gh   h�p���~�  ��u��G;�u�����  _^][��  � �lySS�J�@����P��H  �o\��;Él$�E u����  _^][��  � ���G;É\$��   �  �?Sh�  V���  �L$��Q���   ���  P�L$���  �L$P�G�@�������`  ��  �L$���  ���L?�^\��F�F�D$��\  ��\  ��\  ��\  ��\  �F@  �B�FD  �B�nH�^�^�^�^�n�n �n$�n(�n,�^0�^4�^8�n<�^P�^L�^T�^X�O�ƀ  @;��D$�#����l$�ly�WSS�H��R��H  �wh��;Ét9���   ���8�  ����  ���J�  ��$,  ��P�  V��  U��  ��_^][��  � �����������������HSUV��W�L$ �N�  �N�F\3�3�;���   �  �B�  �?���L?�X\��\  ��\  ��\  ��\  ��\  �@@  �B�hD�HH�8�x�x�X�X�X�X�H�H �H$�H(�H,�X0�X4�X8�H<�XP�XL�XT�XX�  B;Vr���  ��  :�u ��,  �L$ �����,  ��  _^][��H�P�L$��  P�L$@��  P�L$$���  �L$<���  �L$��  ��  �D$ P����  �����   ��W��  ����  ;�t ��,  �L$ �����,  ��  _^][��HË��$   ����  �L$ �t�  _^][��HÐ�������������   S��Uh   ���   h�p�\$3���  ����  VW��p��݃�K�z  3Ɋ��l �$�xl �T$0Rhl4h�p�m �����K  h�p�U�  ���L$ P��  �C3�3���vD3��K\�D$ P��9`  ��  ��u�CF�ǀ  ;�rڍL$ �|�  ��  �C\�v�,����L$ �`�  ��  ����  �D$Ph�4h�p�� ����u�D$�-p!�]�  h�4h�p�� h�4j ���� �����y  ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ�����A  P���  h�   ��\  PQ�} ��ƅ[   �  ���  �T$Rh�4h�p� ����u5�D$��!����Au�D$  �B�D$�uD�ET   ��!�]@��  �D$Ph�4h�p��
 ������  �D$��!����t�D$  �>�L$�MH�|  �D$�|!����Au�D$  �@�L$�MH�W  ���O  ��p<ata<dt6<s�:  �U(�E$R�M PQh�4h�p�5
 �   ���EX�ET�  �U�ERPUh�4h�p�

 ���EP   ��  �M�UQ�ERPh�4h�p��	 ���EL   �  ����  h�4h�p��
 h�4j ����
 P�T�  ������  ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ����u%h�   �M\PQ�	 ��ƅ[   �EP   �,  ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ����uh�   ��\  PR�:	 ����  ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ����uh�   P��\  P�� ���  ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ����u,h�   ��\  PQ� �   ��ƅ[   �EX�ET�0  ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ����u(h�   ��\  PR�> ��ƅ[   �EL   ��   ��4�ϊ��:u��t�Y��:^u������u�3��Ƀ������   h�   P��\  P�� ��ƅ[   �~��tzh�4h�p� h�4j ��� ����tV�x4�ϊ��:u��t�Y��:^u������u�3��Ƀ����u"P���  h�   ��\  PQ�^ ��ƅ[   �\$h   h�p���   �[�  ���R���_^][��   �Ll �h 2h �k ug �i �f Ll  ���������������   SU���D$    �D$    �D$    ��,  �D$$    ��D$     �D$    �D$0    �D$,    �D$(    �D$<    �D$8    �D$4    �  �E��$  j Ph'  ���  �]P�D$�E�D$    ����  VW��4�C����\  �<  ���E`��   �K��t$H�I�����L$H�J�L$L�K��R�I�T$P�����L$T�J�L$X��R�I�T$\�����L$`�J�L$d�K�R�I�T$h�����D$l�J�L$p�   �R�T$t��  �K��$�   �I������$�   �J��$�   ��R�I��$�   ������$�   �J��$�   �K��R�I��$�   ������$�   �J��$�   �K��R�I��$�   ������$�   �J��$�   �   �R��$�   �L  ����   �K��E`Ǆ$�       Ǆ$�       �IǄ$�       �t$x�����L$x�J�L$|�K��R�I��$�   ������$�   �J��$�   ��R�I��$�   ������$�   �J��$�   �   �R��$�   �   ��E`Ǆ$      Ǆ$       �IǄ$�       ��$�   ������$�   �J��$�   �K��R�I��$�   ������$�   �J��$�   �K��R�I��$�   ������$�   �J��$�   �   �R��$�   �ly�|$�HD�D$�T$R�T$PR�Q@�D$�M����P@;��D$�,���_^][���   � �UVW���L$���5  ��,  �(  ��  ���  �L$�l$�I�4ȋEL����\  �H  ���K  �E<�@�GL����!�Z f��E<�WL���@�D���!�< f��E<�OL���@�D���!� f��E@���@�GL����!� f��E@�WL���@�D���!�� f��E@�OL���@�D���!�� f��ED���@�GL����!� f��ED�WL���@�D���!� f��ED�OL���@�D���!�l f��EH���@�GL����!�O f��EH���WL�@�D���!�1 f��mH�  �EH�@�GL����!� f��EH�WL���@�D���!�� f��EH�OL���@�D���!�� f��ED���@�GL����!� f��ED�WL���@�D���!� f��ED�OL���@�D���!�z f��E@���@�GL����!�] f��E@�WL���@�D���!�? f��E@���C  ���K  �E<�@�GL����!� f��E<�WL���@�D���!�� f��E<�OL���@�D���!�� f��E@���@�GL����!� f��E@�WL���@�D���!� f��E@�OL���@�D���!�} f��ED���@�GL����!�` f��ED�WL���@�D���!�B f��ED�OL���@�D���!�$ f��ED���@�GL����!� f��ED���WL�@�D���!��  f��mD�F  �ED�@�GL����!��  f��ED�WL���@�D���!�  f��ED�OL���@�D���!�  f��E@���@�GL����!�n  f��E@�WL���@�D���!�P  f��E@�OL���@�D���!�2  f��E<���@�GL����!�  f��E<�WL���@�D���!���  f��E<���OL�@�D���!���  f��E<���@�GL����!��  f��E<�WL���@�D���!��  f��m<�OL�Dm �D���!��  f�F_^]� ����UW����,  tH�GPhO  ���  �����t1�GS�_PV3���vVSU���t����G��PF;�r�L$j U��  ^[_]� ��������dW���L$T�|$��  �L$@��  ��,  �D$    � �  Vh�� �S�  ���D$����   �ly���   ���R=�� ug�t$�L$0�/�  �ly�T$0RV�H@�Q`���D$0�L$P�M�  �L$0��  �L$Q�L$H��  �L$�m�  �W�L$DRh�  ���  �D$��D$P�+�  ��3��D$�wN�2  ��    ���  +�S��FU�L$�T$�t$�oT���3ۋN����   jh   h�p�����  ��p���3����It��p�   J�< u��@�x�;�r��L$xj h)  ���p�n�  W�L$(�����  �lyP�ˋ��   �R|�L$$��  �D$��t"W�L$<���  P�D$P�L$T�6�  �L$8���  �~���s�  ��F3ۅ�v�Q�����  �F��C;�r�D$�T$�|$ �t$�L$��NI�T$�t$�L$�����][��^t'�lyj�J@�T$DRP�Qd�D$�L$x��j P�Z�  �L$@���  �L$T���  _��d� ���dW���L$T�|$�-�  �L$�$�  ��,  �D$    �@��  Vh�� ���  ���D$����   �ly���   ���R=�� ug�t$�L$0���  �ly�T$0RV�H@�Q`���D$0�L$DP���  �L$0�$�  �L$DQ�L$ �&�  �L$D��  �W�L$Rh�  �k�  �D$��D$P���  ��3��D$�wN��   ��    ���  +�S��FU�L$�T$�t$�_X���N��tq�L$xj h)  �Y�  �ly��V�ˋ��   �P|�D$��t�L$VQ�L$,�>�  �~����  ��F3ۅ�v���R���  �F��C;�r�D$�|$ �T$�t$�L$��NI�T$�t$�L$�b���][��^t'�lyj�Q@�L$QP�Rd�T$�L$x��j R�k�  �L$���  �L$T���  _��d� ����h  SUV��W�L$�t$$�7�  h 5�L$@���  P��  ���L$<��  �nM�l$,��  �Dm �|� ���|$(��|$(��$|  �X�  �L$$���D$0    y\��t_��`  �ly�΋��   �PxS����  ��u�ly���   ���R(����u��#�ly�΋��   �R=G  u^���D$0   u&��  �����1  �ly�΋��   ��`  P�R|�L$$��,  ��t6�GP��u/�lyj j V�BT�P4��   �D$$�Hl��   �Ph�4��  �lyj V�QT�R,���荄$   ��P�f�  P�L$�l�  ��$   �P�  ��\$d�G�\$h�G�L$dQh�  �\$t�L$���  h  �?h�  �L$��  �O\�G\��tHP��$�   �O�  Ph�  �L$���  ��$�   �d�  jh�  �L$�D�  jh�  �L$�4�  �T$��R��  �lyjj V�HT�Q4�G�� ������@��   �WH�L$4R��  �lyjV�HT�Q,���荔$�   ��R�b�  P�L$�h�  ��$�   �L�  �G�L$Ph�  ���  �L$Q���~�  �T$4j �D$PRP�L$|�D$X�  �D$\    �D$`    ��  P�����  �L$p�0�  �lyjjV�QT�R4���L$4�C�  ��lyj jV�HT�Q4���GL���  �G�� ����@t$�G�� ����@t�G�� ����@��   �lyjV�QT�R,���荄$P  ��P�\�  P�L$�b�  ��$P  �F�  �G�\$X�G�\$\�G�L$XQh�  �\$h�L$���  h  �?h�  �L$��  ��\  ��\  ��tHP��$�   �>�  Ph�  �L$��  ��$�   �S�  jh�  �L$�3�  jh�  �L$�#�  �T$��R���  �lyjjV�HT�Q4��lyj jV�BT�P4�GT�ly���QT��tOjV�R,���荄$(  ��P�W�  P�L$�]�  ��$(  �A�  �L$Q����  �lyjjV�BT�P4�j jV�R4�GX�����  �G �� ����@t$�G$�� ����@t�G(�� ����@��   �lyj	V�BT�P,����$�   ��Q����  P�L$��  ��$�   ��  �G �\$<�G$�\$@�G(�T$<�L$Rh�  �\$L�'�  h  �?h�  �L$���  ��\  ��\  ��tBP�L$|��  Ph�  �L$��  �L$x��  jh�  �L$��  jh�  �L$��  �D$��P�V�  �lyjj	V�QT�R4��lyj j	V�HT�Q4��\  �ly��\  �����BT��   jV�P,����$  ��Q����  P�L$��  ��$  ��  S��$�   ���  Ph�  �L$�G�  ��$�   ���  jh�  �L$���  �T$��R��  �lyjjV�HT�Q4�j jV�P4��\  �ly���QT��twjV�R,���荄$<  ��P��  P�L$��  ��$<  ��  S��$�   �2�  Ph�  �L$��  ��$�   �G�  �L$Q����  �lyjjV�BT�P4�j jV�R4��\  ��\  �����ly�HTtwjV�Q,������$d  ��R�k�  P�L$�q�  ��$d  �U�  S��$�   ��  Ph�  �L$�	�  ��$�   ��  �D$��P�q�  �lyjjV�QT�R4�j jV�Q4�D$<����u��$|  j j V���  jj���o�  �T$$�L$,��Bh�4��L$(M��  �l$,��L$(�<����L$諾  _^][��h  � ����������������DW���L$�|$���  ��,  �u�L$�k�  _��D� �D$LSUVP�������GH��   �@����@�L$X�D$�w\�p  ��te�L$\j h)  ���  �ly��`  ��Q���   ���P|��x  ����  �苆p  3ۅ�v���R�{�  ��p  ��C;�r�|$�L$X�D$��  H�L$X�D$�s����_K��   �[�,�����|$�w\�L$\j h�  ��>�  �L$,����  �ly�D$,PW�Q@�R`���L$,Q�L$D��  �L$,�G�  �T$@�L$R�I�  �L$@�0�  ��`  �L$Vh�  ��  jh�  �L$ �{�  �ly�T$jR�H@W�Qd�D$���Hh����R�3�  K��  ���=����L$�˼  ^][_��D� ���8S��W�\$�C�PQ�9�  �������|$u(h�5�L$4���  P�(�  ���L$0���  _[��8� �T$HUVR�L$<��  �lyP���   ���R|�L$8���  �lyj h�  W�HH�Q|�ly�D$8j h�  �BHW�P|�����L$8�t$0h�5�W�  P���  ���L$8�u�  �K�CP���D$     v}���΋P0����\  u/��t��p�X�h��P�p�X�(����w�_�\$�o�!��t�P�0���p�x��u �}�U�U�T$ �s�|$��PB��;։T$ r���CH3Ʌ�v)�T$,������A�.���/�n�o�v�w�3;�rߋ|$��X  ��t(h�5�L$<�j�  P���  ���L$8��  W��������P  ��t(hl5�L$<�8�  P���  ���L$8�V�  W��������L  ��t(hT5�L$<��  P��  ���L$8�$�  W���|�����T  ��t-h 5�L$<���  P�^�  ���L$8���  �L$LWQ���������`  ��t(h<5�L$<��  P�'�  ���L$8��  W��������d  ���M  �C ���B  ���3�  ����  ���D$4�(  �lyj j�ϋ��   �P�K 3��ɉD$ ��  �spP�Kt�.�  3�;���  �h3�;�v�hA�T���h;�r�H�T$P;ʉT$�  �P�|$�,��y��L$�l$$;�u�:�|$�
�L��L$���H3҅���   �H�L$(��|$�L$(�\$0�	��ˋ;�u9ytE9iu9ytF�y�l$$;�u;\$tD�I�l$$;�t
;�u;|$t>�|$(�HB��;щ|$(r��O�H�����+�H����   ��H����   ��H����   ��H�����B��L$PA�L$P�\$�|$�HG�׉|$;�������|$�T$P�H;�ud�N�����    3҉�h3Ʌ�v(�h�|�  u�h���l� ����   @B�.�hA;�r؋L$,�@Q�L$4�Q�KpPj Q�L$Hj ��  �$h5�L$<�[�  �T$8R�q�  ���L$8�u�  �D$ �K @;��D$ �����L$4�8�  �t$Ljj j W�����  j h�  ���x�  h¸�?jj���x�  �lyj j�ϋ��   �Rj W�����  ^]_[��8� ���D$ S�\$4��UV�t$@3�W�zp���T$vO��T$�D$,�jP3ҋ ����ŋk��v�k�l� ;hu�n�L� �kB;�r�l$,�D$0��A;ȉl$,r��K3��N�S�ɉVv�L$4�S�n��@���T���V;�r�N3�3�;�v�N@�T���N;�r�F�T$,;T$4�  �NH;Ћ,��l$Du�	�L$0�
�T��T$0�ʋF3҅���   �F�D$@��L$0�D$@�\$8� ��Ë;�u9HtE9hu9HtQ�H�l$D;�u;\$0tO�@�l$D;�t
;�u;L$0tU�L$@�FB��;ЉL$@r��f�F������F�����B�F����   �(�F������   �O��F����F����   ��N�����A��D$,@�D$,�T$4�FB;ЉT$4������T$,�F;�un�_�����    3ɉ�V3���v&�V�<� u�V��������   @A��V@;�rڋD$<�T$8P�F��L$RP�Qp�L$4j Rj ��  _^][���  h5�L$�i�  �D$P��  ���L$��  _^][���  �����������,  SU��V3�W�L$|�l$d�U�  ��,  �l$4� �l$ �l$$�l$u��$D  ��$@  PQ���������  �ly�UU�B��Q��H  �ly��D$$U�BU��Q��H  �ly�K�D$LU�BU��Q��H  �ly�K�D$DU�BU��Q��H  �D$T��T  ��0;�t��,  �t��$@  ��R�<���h�5��$�  �K�  P���  ����$�  �f�  �C�sT;ŉt$�l$H��  ��$�   �D�  �L$h�;�  9nu!���L$h�t$観  ��$�   蚳  �  jh   h�p���R�  ��p���3����It��p�   J�< u��@�p�;�r��|$����p�GPQ�и  �������t$,��  U��$�  �r�  �lyP�΋��   �R|��$�  ��  �lyj h�  V�HH�Q|�ly�D$`j h�  �BHV�P|��`  �D$t3���;ȉD$@t ��,  t�OQhO  �;�  ���D$@3���X  �D$P;�t ��,  t�WPRh'  ���j�  �D$P3���L  �D$(;ȉD$`�d  j h)  ����  U��$0  ����  �lyP���   ���R|��$,  ��  ���<�  h�� �D$d�~�  ���D$(���  �ly���   ���R=�� ��   �|$(��$�  �S�  �ly��$�  RW�H@�Q`����$�  ��$  P�h�  ��$�  蜱  ��$  Q��$�   蘱  ��$  �|�  jh�  ��$�   �ٳ  U��$�  ��  Ph�  ��$�   ��  ��$�  ��  �ly��$�   jQ�B@�T$0R�Pd�D$4��3���WP葵  ��L$(Q��  ��3��|$(�3���D$4��WRP�G�  �K�T$,��WQR�5�  �C�L$<��WPQ�#�  �D$@��$�|$<�|$L�H�P;ω|$�T$D�|$�  �D$\�D$8�  �D$0�L$`��t
�T$R��  �D$D�KP�D$X    �(�l� ���EL��vp�t$<�T$T�E�v����|$4���<9 u=�|$�4��sH�I����9�>�y�~�I�N�t$<��|$4F���t$<��   �L$X�}LA��;ωL$Xr��EL����\  uL��t-�U�D$�u$�}(���U �4������|$0��W�w�G�S�M(�D$�U$�u ���}���4��х�t�M$�D$�U����M�D$�U$���u �����t$0��F�N�N�D$@��t�L$QUP���o����D$P���z  �ELǄ$�       ����\  Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       �d  ���C`��   �M,��$  �I������$  �Q��$  �I��$  �M0�I������$  �Q��$  �I��$  �M4�I������$  �Q��$   �I��$$  �M8�I�����$(  �   �P��$,  �@��$0  �  �M8��$d  �I������$d  �J��$h  �M4�R�I��$l  ������$p  �J��$t  �M0�R�I��$x  ������$|  �J��$�  �M,�R�I��$�  ������$�  �J��$�  �   �R��$�  �W  ����   �M,�C`Ǆ$       Ǆ$�       �IǄ$�       ��$�   ������$�   �J��$�   �M0�R�I��$�   ������$�   �J��$�   �M4�R�I��$�   ������$�   �J��$�   �   �R��$�   �   �M4�C`Ǆ$`      Ǆ$\      �IǄ$X      ��$4  ������$4  �J��$8  �M0�R�I��$<  ������$@  �J��$D  �M,�R�I��$H  ������$L  �J��$P  �   �R��$T  �ly��$�   �HD�D$��$�   R�T$TPR�Q@����P  ���L  ��,  @�?  �E�L$ �<� �  �L$,��    +ЋCXj h)  �<��.�  ������   �lyW���   ���R|���k�  �M�T$ ���D$����   h�� 蛮  ���D$����   �ly���   ���R=�� ��  �t$��$�  �p�  �ly��$�  RV�H@�Q`����$�  ��$  P腪  ��$�  蹪  ��$  Q�L$l踪  ��$  蜪  �D$��t�t$8WV�L$p�U�  �L$LAF�L$L�t$8�E�L$ ����t
�T$R���  ��T  ���H  ��,  ��;  �E�L$$�<� �  �{\�L$,�@j h)  �4�����ծ  ������   �ly��`  V�ϋ��   �R|����  �M�T$$j h�  ���L$4蓮  ��$�  ���E�  �ly��$�  RW�H@�Q`����$�  ��$�  P�Z�  ��$�  莩  ��$�  Q��$�   芩  ��$�  �n�  Vh�  ��$�   �,�  jh�  ��$�   蹫  �ly�L$|jQ�B@W�Pd�U�Ch����Q���q�  �U�D$$����t
�T$R��  �l$D�L$�D$�t$0�Q��@��;l$D�D$�t$0�Q����D$��t=�T$L�L$hRh�  �0�  �ly�T$hjR�H@�D$P�Qd�L$ ��j Q�L$4��  �D$@��t*�t$,j P��� �  ��T$R�T�  ���D$    ������t$,�l$�D$<�΋URP�l�  ��d  ����   �C ����   ���L�  ���%�  ���D$8��   �lyj j���   ���R�C �D$    ��vg�D$�KtP�H�  �L$��Q���   �6�  ��tD��t@�T$H�O;�u%�L$\�T$P�D$XWP�EQ�MR�T$LPQR�������D$�K @;��D$r��|$8����  j��誼  �D$d��$@  jPj V����  j h�  ����  h¸�?jj����  �lyj j���   ���Rj V����  ���L$h�t$d�l$��  ��$�   ��  ��3�D$H�K@;��D$H�����D$$P��  �L$$Q�	�  �T$<R���  �D$$P���  ���L$|蹦  _^][��,  � h�5��$�  ��  P�5�  ����$�  ��  �L$h�}�  ��$�   �q�  뭐����������������,  SU��V3�W�L$|�l$d�ť  ��,  �l$4�@�l$ �l$$�l$u��$D  ��$@  PQ���T�����  �ly�UU�B��Q��H  �ly��D$$U�BU��Q��H  �ly�K�D$LU�BU��Q��H  �ly�K�D$DU�BU��Q��H  �D$T��T  ��0;�t��,  �t��$@  ��R����h�5��$�  軻  P�E�  ����$�  �ֻ  �C�sX;ŉt$�l$H��  ��$�   贤  �L$h諤  9nu!���L$h�t$��  ��$�   �
�  �  jh   h�p���¼  ��p���3����It��p�   J�< u��@�p�;�r��|$����p�GPQ�@�  �������t$,��  U��$�  ��  �lyP�΋��   �R|��$�  ���  �lyj h�  V�HH�Q|�ly�D$`j h�  �BHV�P|��`  �D$t3���;ȉD$@t ��,  t�OQhO  諧  ���D$@3���X  �D$P;�t ��,  t�WPRh'  ���ڨ  �D$P3���P  �D$(;ȉD$`�X  j h)  ��耨  U��$0  ����  �lyP���   ���R|��$,  ��  ��謦  h�� �D$d��  ���D$(����   �ly���   ���R=�� ��   �|$(��$�  �â  �ly��$�  RW�H@�Q`����$�  ��$  P�آ  ��$�  ��  ��$  Q�L$l��  ��$  ��  jh�  �L$p�O�  U��$�  �"�  Ph�  �L$p蓥  ��$�  �7�  �ly�L$hjQ�B@�T$0R�Pd�D$4��3���WP��  ��L$(Q�a�  ��3��|$(�3���D$4��WRP�ô  �K�T$,��WQR豴  �C�L$<��WPQ蟴  �D$@��$�|$<�|$L�H�P;ω|$�T$D�|$�  �D$\�D$8�  �D$0�L$`��t
�T$R蔾  �D$D�KP�D$X    �(�l� ���EL��vp�t$<�T$T�E�v����|$4���<9 u=�|$�4��sH�I����9�>�y�~�I�N�t$<��|$4F���t$<��   �L$X�}LA��;ωL$Xr��EL����\  uL��t-�U�D$�u$�}(���U �4������|$0��W�w�G�S�M(�D$�U$�u ���}���4��х�t�M$�D$�U����M�D$�U$���u �����t$0��F�N�N�D$@��t�L$QUP��������D$P���z  �ELǄ$�       ����\  Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       �d  ���C`��   �M,��$  �I������$  �Q��$  �I��$  �M0�I������$  �Q��$  �I��$  �M4�I������$  �Q��$   �I��$$  �M8�I�����$(  �   �P��$,  �@��$0  �  �M8��$d  �I������$d  �J��$h  �M4�R�I��$l  ������$p  �J��$t  �M0�R�I��$x  ������$|  �J��$�  �M,�R�I��$�  ������$�  �J��$�  �   �R��$�  �W  ����   �M,�C`Ǆ$       Ǆ$�       �IǄ$�       ��$�   ������$�   �J��$�   �M0�R�I��$�   ������$�   �J��$�   �M4�R�I��$�   ������$�   �J��$�   �   �R��$�   �   �M4�C`Ǆ$`      Ǆ$\      �IǄ$X      ��$4  ������$4  �J��$8  �M0�R�I��$<  ������$@  �J��$D  �M,�R�I��$H  ������$L  �J��$P  �   �R��$T  �ly��$�   �HD�D$��$�   R�T$TPR�Q@����L  ���R  ��,   �E  �E�L$ �<� �  �L$,��    +ЋCTj h)  �<�誡  ������   �lyW���   ���R|����  �M�T$ ���D$����   h�� ��  ���D$����   �ly���   ���R=�� ��  �t$��$�  ��  �ly��$�  RV�H@�Q`����$�  ��$  P��  ��$�  �5�  ��$  Q��$�   �1�  ��$  ��  �D$��t �t$8WV��$�   �˞  �L$LAF�L$L�t$8�E�L$ ����t
�T$R�u�  ��T  ���H  ��,  ��;  �E�L$$�<� �  �{\�L$,�@j h)  �4�����K�  ������   �ly��`  V�ϋ��   �R|��胞  �M�T$$j h�  ���L$4�	�  ��$�  ��軚  �ly��$�  RW�H@�Q`����$�  ��$�  P�К  ��$�  ��  ��$�  Q��$�   � �  ��$�  ��  Vh�  ��$�   袝  jh�  ��$�   �/�  �ly�L$|jQ�B@W�Pd�U�Ch����Q����  �U�D$$����t
�T$R��  �l$D�L$�D$�t$0�Q��@��;l$D�D$�t$0�K����D$��tC�T$L��$�   Rh�  補  �ly��$�   jR�H@�D$P�Qd�L$ ��j Q�L$4膞  �D$@��t*�t$,j P���p�  ��T$R�ğ  ���D$    ������t$,�l$�D$<�΋URP�ܞ  ��d  ����   �C ����   ��輟  ��蕟  ���D$8��   �lyj j���   ���R�C �D$    ��vg�D$�KtP踑  �L$��Q���   覑  ��tD��t@�T$H�O;�u%�L$\�T$P�D$XWP�EQ�MR�T$LPQR�������D$�K @;��D$r��|$8���S�  j����  �D$d��$@  jPj V����  j h�  ��脝  h¸�?jj��脜  �lyj j���   ���Rj V����  ���L$h�t$d�l$聘  ��$�   �u�  ��3�D$H�K@;��D$H�����D$$P胪  �L$$Q�y�  �T$<R�o�  �D$$P�e�  ���L$|�)�  _^][��,  � h�5��$�  �[�  P襩  ����$�  �v�  �L$h��  ��$�   ��  뭐����������������L  SU��V3�W�L$x�l$t�5�  ��,  �l$D���l$(�l$,�l$u��$d  ��$`  PQ��������  �ly�UU�B��Q��H  �ly��D$(U�BU��Q��H  �ly�K�D$\U�BU��Q��H  �ly�K�D$LU�BU��Q��H  �D$\��T  ��0;�t��,  �t��$`  ��R����h�5��$�  �+�  P赯  ����$�  �F�  �K�C\;͉l$H��  ��x  ��p  `  �L$8�T$�D$<��  ��$�   ��  ��$�   ���  �D$9(u9�T$<�ȋD$8�։L$ƍ�$�   �T$<�D$8�J�  ��$�   �>�  �  �L$<jh   h�p���  ��p���3����It��p�   J�< u��@�p�;�r��|$����p�QR�s�  �������t$4�	  U��$�  ��  �lyP���   ���R|��$�  �'�  �lyj h�  V�HH�Q|�ly�D$tj h�  �BHV�P|��$�   ��`  ���D$P    ��t��,  t�QhO  �ژ  ���D$P��X  �D$L    ��t��,  t�j Rh'  ����  �D$L��T  �D$p    ���  j h)  ��诙  U��$P  ���0�  �lyP���   ���R|��$L  �B�  ���ۗ  j h�  �ΉD$x�i�  ������   ��$�  ��  �ly��$�  RV�H@�Q`����$�  ��$  P�(�  ��$�  �\�  ��$  Q�L$|�[�  ��$  �?�  �T$<�L$xRh�  ���  jh�  ��$�   艖  �ly�T$xjR�H@V�Qd�Ch�L$T������R�A�  ��L$D3���WPQ�>�  �S�D$4��WRP�,�  �K�T$D��WQR��  �D$\�T$4��$�|$X��;ǉ|$T�|$\�|$�|$�L$`�|$$��  ��  �D$@�D$d�D$l�D$0�L$p��t
�T$$R� �  �D$`�KP�D$     �(�l� ���EL��vl�T$h��E����t$D���<1 u=�t$�<1��sH�I����9�>�y�~�|$X�IG�N��t$D�|$X����   �L$ �uLA��;ΉL$ r��EL����\  uz��t;�D$�u$�U�4����U ��$D  �u(�����t$0���$D  �V�N�F�s�D$�u �U(�4����U$��$�  �u�����t$0���$�  �V�N�F�8��t�U$�D$���U��M�D$�U$���u �����t$0��F�N�N�D$P��t�L$$QUP���-����D$L���~  �ELǄ$�       ����\  Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       Ǆ$�       �d  ���C`��   �M,��$  �I������$  �Q��$  �I��$  �M0�I������$   �Q��$$  �I��$(  �M4�I������$,  �Q��$0  �I��$4  �M8�I�����$8  �   �P��$<  �@��$@  �  �M8��$t  �I������$t  �J��$x  �M4�R�I��$|  ������$�  �J��$�  �M0�R�I��$�  ������$�  �J��$�  �M,�R�I��$�  ������$�  �J��$�  �   �R��$�  �W  ����   �M,�C`Ǆ$p      Ǆ$l      �IǄ$h      ��$D  ������$D  �J��$H  �M0�R�I��$L  ������$P  �J��$T  �M4�R�I��$X  ������$\  �J��$`  �   �R��$d  �   �M4�C`Ǆ$      Ǆ$      �IǄ$      ��$�   ������$�   �J��$�   �M0�R�I��$�   ������$�   �J��$�   �M,�R�I��$�   ������$�   �J��$   �   �R��$  �ly��$�   �HD�D$$��$�   R�T$PPR�Q@�|$d����L  ���^  ��,   �Q  �E�L$(�<� �(  ��    j +ЋCTh)  ���L$(�L$<��  ������   �ly�L$ Q�΋��   �P|����  �U�L$(���D$����   h�� �M�  ���D$����   �ly�ȋ��   �R=�� ��  �t$��$�  �"�  �ly��$�  RV�H@�Q`����$�  ��$   P�7�  ��$�  �k�  ��$   Q��$�   �g�  ��$   �K�  �D$��t$�D$ �t$dPV��$�   ���  �L$TAF�L$T�t$d�M�T$(����t
�D$$P觩  ��P  ����  ��,  @��  �E�L$,�<� �[  ��    j +ЋCXh)  ���L$(�L$<�x�  �����.  �ly�L$ Q�΋��   �P|��豏  �U�L$,���D$����   h�� ��  ���D$����   �ly�ȋ��   �R=�� ��   �t$��$�  趋  �ly��$�  RV�H@�Q`����$�  ��$(  P�ˋ  ��$�  ���  ��$(  Q��$�   ���  ��$(  �ߋ  �1�T$R賑  ���D$    �����T$R虑  ���D$    �,�D$��t$�D$ �t$@PV��$�   �^�  �L$\AF�L$\�t$@�M�T$,����t
�D$$P��  �D$`�L$�t$0����D$`�D$$��@�t$0;D$$������D$��tC�T$T��$�   Rh�  荍  �ly��$�   jR�H@�D$ P�Qd�L$$��j Q�L$<�p�  �D$��tC�T$\��$�   Rh�  �B�  �ly��$�   jR�H@�D$P�Qd�L$ ��j Q�L$<�%�  �D$P��t�t$4j P����  ��t$4�T$�΋PW蚏  ��d  ����   �C ����   ���z�  ���S�  ���D$@��   �lyj j���   ���R�C 3��v\U�Kt耂  U���   ���r�  ��tA��t=�L$H�;�u+�T$h�L$P�D$pWR�T$PQ�L$L��P�D$XRP���U����C E;�r��|$@���"�  j����  �L$t��$`  jQj V���ѫ  j h�  ���S�  h¸�?jj���S�  �lyj j�΋��   �Pj V���ԫ  �L$8�T$��  �t$t�t$<��ЉL$8��$�   �t$<�T$�1�  ��$�   �%�  ��  3�D$H�K@;��D$H�x����L$,Q�0�  �T$,R�&�  �D$LP��  �L$(Q��  ���L$x�ֈ  _^][��L  � h�5��$�  ��  P�R�  ����$�  �#�  ��$�   藈  ��$�   苈  몐��������S��VW�KP�{  �Kd�w  �Kt�w  ���  �x�  3��   ���  ���   ���   ���   ���   ���   ���   �C�C ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ��  ��  ��  ��$  �6������  ���  ��   ��  ��  ��  ��  ǃ�     ǃ�  �  �C4�C8�C<�C@�CD�C,�C0�CH�CL���  ���  ���+����  ���������ȋÃ��_^[Ð�����SV��W�^P����}  ����  ���  ���  ��t	W��  �����  �    萤  �Nt�w  �Nd�w  ���z  _^[Ð����S��U�C@�k@��tK�CW3���v0V3��E ��x  ��x  ��t	P�ʘ  ���CG�ƀ  ;�r�^U貘  ���E     _][Ð���S��U�C8�k8��tB�CW3���v'V3��E �L�D��t	P�p�  ���CG��;�r�^U�[�  ���E     _][Ð������������S��U�C<�k<��tB�CW3���v'V3��E �L�D��t	P��  ���CG��;�r�^U���  ���E     _][Ð������������UW���GL�oL��tf�O S3ۅ�vDV�p�N��F���t	P贗  ���> t	V覗  ���N�F��t	P蓗  ���G �� C;�r�^U�~�  ���E     �G     [_]Ð��������VW���w������������������B����F4�~4��t	W�2�  ���F,�    �~,��t	W��  ���F0�    �~0��t	W� �  ���FD�    �~D��t	W��  ���FH��H���    t	V�Ζ  ���    _^Ð�UVW��3�GL;��b  �t$���9.�Q  S�_dhD6����t  ���  �FI���  �$�<� ;ŉl$�  �,������F���   �(�D�NP���   �)�L�VQ���   �*�T���  Rh46P謵  �����  ��P�[t  �D$�N@��;��D$r��  ;���  �F���   ���D�NP���   ���L�VQ���   ���T���  Rh46P�7�  �����  ��P��s  �FE;�r��*  ;ŉl$�  �,������F���   �(�D�NP���   �)�L���  Qh(6P�Ӵ  �����  ��P�s  �D$�N@��;��D$r��  ;���  �V���   ���T�FR���   ���DP���  h(6P�o�  �����  ��P�s  �FE;�r��b  ;ŉl$�V  �,������N���   �)�L�VQ���   �*�T���  Rh6P��  �����  ��P�r  �D$�N@��;��D$r���   ;���   �F���   ���D�NP���   ���L���  Qh6P觳  �����  ��P�Vr  �FE;�r��   ;ŉl$��   �,������V���   �*�T���  Rh6P�T�  �����  ��P�r  �D$�N@��;��D$r��?;�v;�F���   ���DP���  h6P��  �����  ��P�q  �FE;�r�hP4���q  �   [_^]� ��� �� �� f� �� .� �� � ����SUV��W���  H���~  �$�� �D$�N0�~H�n$���   ���   ������l$���   �DP��DP�D$� �D(P�A�DP�G�DP�D$(�@�D(P�A�I�DP�G�T�DP�D$4�@�D(P�GR�T$<�L�BQ�   �D$�N0�~H�n$���   ���   �����A�l$���   �DP�G�DP�D$�@�D(P�A�DP�G�DP�D$(�@�D(P�A�	�DP�G�T
�DP�D$4�@�D(P�R�T$<�L�Q�L(���  Qh�6R�P�  ��8�,  �D$�NH���   �~$���ǋ��   ��\S��\S�Y�\S�X�\;S�Y�I�\S�X�@�T�\;S�L8RQ���  h�6R�ܰ  ��(�  �D$�NH���   �~$���ǋ��   �Y�\S�X�\;S�Y�\S�X�\;S�Y�	�\S�X� �T
�\;S�LRQ���  h�6R�h�  ��(�D  �D$�N0���   �~$���ǋ��   ��\S��\S�Y�\S�X�\;S�Y�I�\S�X�@�T�\;SR�L8�Z�D$�N0���   �~$���ǋ��   �Y�\S�X�\;S�Y�\S�X�\;S�Y�	�\S�X� �T
�\;SR�LQ���  h\6R蘯  ��(�w�D$�N$������   ��TR�P�T
R�P�@�T
R�L�0�D$�N$������   �P�T
R�P�T
R�P� �T
R�LQ���  hH6R��  �����  �NdP��m  _^][� ��}� � �� <� �� � }� �� ����SUV��W���  H����  �$�H� �D$�N0�~H�n$���   ���   ������l$���   �DP��DP�D$� �D(P�A�I�DP�G�T�DP�D$(�@�D(P�GR�T$0�L�BQ�x�D$�N0�~H�n$���   ���   �����A�l$���   �DP�G�DP�D$�@�D(P�A�	�DP�G�T
�DP�D$(�@�D(P�R�T$0�L�Q�L(���  Qh(7R軭  ��,��  �D$�NH���   �~$���ǋ��   ��\S��\;S�Y�I�\S�X�@�T�\;S�L8RQ���  h7R�W�  �� �p  �D$�NH���   �~$���ǋ��   �Y�\S�X�\;S�Y�	�\S�X� �T
�\;S�L8RQ���  h7R��  �� �  �D$�N0���   �~$���ǋ��   ��\S��\;S�Y�I�\S�X�@�T�\;SR�F�D$�N0���   �~$���ǋ��   �Y�\S�X�\;S�Y�	�\S�X� �T
�\;SR�L8���  Qh�6R�G�  �� �c�D$�N$������   ��T
R�P�@�T
R�$�D$�N$������   �P�T
R�P� �T
R�L���  Qh�6R��  �����  �NdP�j  _^][� �M� �� ]� �� %� m� �� �� ����������<  SUVW��3�� }  h�7�L$@�|$�\$$����  P菒  ���L$<�#�  �N�F@;ω|$�   ��p  �L$�3��҉D$��  �Q���V4�<�������tp�FL��ti�W���< t]���   G�ǉ��   �?��  ���  ��  ���   �D$43��L$$�D$8�D$(�l$4�t$$��!��  P跑  ���I  ���  ����   ��  ����   ���   ��   �G;���   ��    +ЋF8��觏  ����   �Gj�L$Ph   ��    Q+ЋF8���L�  �L$LQ�v  �O����t-��$T  ��t"��  ��tP���  Qh|7U� �  ������  Pht7U��  ��U�Nd�h  ���  ��tv���  @tm�G;�tf��    +ЋF<����  ��tN�Gj�L$Ph   ��    Q+ЋF<��蘏  �L$LQ��u  �����  Phl7U�i�  ���NdU�h  ���  ��tZ�G�L$ ;�tOj�T$P�@h   R���F@����`  �4�  �L$LQ�ju  �����  Ph`7U��  ���NdU�g  ��W�o�_���T$ t�G��P������Lu�OQ��������W��R��������   B���   �?u=���  t4���   �D$,3��L$<�D$0�D$@�l$,�t$<��!觪  P�m�  ���D$�L$�D$�@;D$�����D$�V���  @;L$�D$������T$���  RhP7W��  ���NdW��f  _^][��<  � ����<  SUVW��3�� }  h�7�L$@�|$�\$$���e�  P��  ���L$<背  �N�F8;ω|$�  �H�L$�3��҉D$��  �Q���V4�<�������tp�FL��ti�W���< t]���   G�ǉ��   �?��  ���  ��  ���   �D$43��L$$�D$8�D$(�l$4�t$$��!�T�  P��  ���I  ���  ����   ��  ����   ���   ��   �G;���   ��    +ЋF8���
�  ����   �Gj�L$Ph   ��    Q+ЋF8��诌  �L$LQ��r  �O����t-��$T  ��t"��  ��tP���  Qh|7U�c�  ������  Pht7U�L�  ��U�Nd� e  ���  ��tv���  @tm�G;�tf��    +ЋF<���R�  ��tN�Gj�L$Ph   ��    Q+ЋF<�����  �L$LQ�1r  �����  Phl7U�̥  ���NdU�d  ���  ��tZ�G�L$ ;�tOj�T$P�@h   R���F@����`  藋  �L$LQ��q  �����  Ph`7U�h�  ���NdU�d  ��W�o�_���T$ t�G��P�������Lu�OQ���z�����W��R�=������   B���   �?u=���  t4���   �D$,3��L$<�D$0�D$@�l$,�t$<��!�
�  P�Ћ  ���D$�L$�D$�@;D$�����D$�V��@;L$�D$������T$���  RhP7W聤  ���NdW�5c  _^][��<  � ����������<  SUVW��3�� }  h�7�L$@�|$�\$$���ň  P�O�  ���L$<��  �N�F<;ω|$�  �H�L$�3��҉D$��  �Q���V4�<�������tp�FL��ti�W���< t]���   G�ǉ��   �?��  ���  ��  ���   �D$43��L$$�D$8�D$(�l$4�t$$��!败  P�z�  ���I  ���  ����   ��  ����   ���   ��   �G;���   ��    +ЋF8���j�  ����   �Gj�L$Ph   ��    Q+ЋF8����  �L$LQ�Eo  �O����t-��$T  ��t"��  ��tP���  Qh|7U�â  ������  Pht7U謢  ��U�Nd�`a  ���  ��tv���  @tm�G;�tf��    +ЋF<��貇  ��tN�Gj�L$Ph   ��    Q+ЋF<���[�  �L$LQ�n  �����  Phl7U�,�  ���NdU��`  ���  ��tZ�G�L$ ;�tOj�T$P�@h   R���F@����`  ���  �L$LQ�-n  �����  Ph`7U�ȡ  ���NdU�|`  ��W�o�_���T$ t�G��P�M�����Lu�OQ���������W��R�������   B���   �?u=���  t4���   �D$,3��L$<�D$0�D$@�l$,�t$<��!�j�  P�0�  ���D$�L$�D$�@;D$�����D$�V��@;L$�D$������T$���  RhP7W��  ���NdW�_  _^][��<  � ����������4  SUV��W� }  h�7�L$8�D$    �\$���#�  P譇  ���L$4�A�  �F�~43�;��L$��  �3ɋ��tk�FL;�td�W��9tY���   @�?���   ��  ���  �|  �D$���   �L$ �D$,�l$�L$0�t$,��!�9�  P���  ���E  9��  ��   9�  ��   ���   ��   �G;���   �V8��    +ȍ���  ����   j�D$H�V8h   P�G��    +ȍ�蘅  �D$DP��k  �O����t-��$L  ��t"��  ��tP���  Qh|7U�L�  ������  Pht7U�5�  ��U�Nd��]  ���  ��tv���  @tm�G;�tf�V<��    +ȍ��;�  ��tNj�D$H�V<h   P�G��    +ȍ���  �D$DP�k  �����  Phl7U赞  ���NdU�i]  ���  ��tZ�G�L$;�tO�@j�L$Hh   ��Q�N@����`  耄  �T$DR�j  �����  Ph`7U�Q�  ���NdU�]  �G�o�_�D$���t�OQ���������Lu�W��R�c�����G��P�&������   B���   �?u=���  t4���   �D$$3��L$4�D$(�D$8�l$$�t$4��!��  P蹄  ���D$�D$�N��P@;��D$�0����T$���  RhP7W腝  ���NdW�9\  _^][��4  � ������������V���  ��t_�FH��tX���  ��t,�F0��t%���  ��tǆ�     �   ǆ�     �u���  ��tǆ�     �_ǆ�     �S���  ��t)�F0��t"���  ��tǆ�     �,ǆ�     � ���  ��tǆ�     �
ǆ�     ��$  W�|$�FL    ��t��   ��tW����s����u��   ��   ��t�D$��PW�����?��  ��t�L$QW���?����&��  ��t�T$��RW�������D$��PW�W����Nd�oZ  ���  _��t���=����   ^� ������xV��W�F���;�v��3��@�~H�lyWW�Q��P��H  ��;ǉFDuh<8�*h  ��3�_^��x� �ly�FWW�Q��P��H  ��;ǉFHuh08��g  ��3�_^��x� �NQ�Km  ��;ǉD$uh$8��g  ��3�_^��x� ��$�   PR���8����u!h8�g  �D$P�1o  ��3�_^��x� �FSU3�;ǉl$�}  �ly�D$`    �D$\    �D$X    �D$l    �D$h    �D$d    �D$x    �D$t    �D$p    Ǆ$�       Ǆ$�       �D$|    �QD�L$�D$XPUQ�R<���  ����t6�D$X�-p!�D$d�-p!�\$(�D$p�-p!�\$4�D$|�-p!�\$@��T$d�D$p�L$|�T$(�D$X�D$4�L$@���  ��t%�T$\�D$h�L$t�T$P��$�   �D$,�L$8�T$D�;�D$\�-p!�\$P�D$h�-p!�\$,�D$t�-p!�\$8ل$�   �-p!�\$D�F$ǋX�H���   +����3҃�3Ƀ�;��_  �ÉT$���D$ �l$�FD���u@�E ������!����t,�E�d$P����!����t�FH���8���   H���   ��uC�E �d$(����!����t-�E�d$,����!����t�FH���T8���   H���   ��uC�E �d$4����!����t-�E�d$8����!����t�FH���T8���   H���   �D$ ��tH��uC�E �d$@����!����t-�E�d$D����!����t�FH���T8���   H���   ��+�t�l$���   B��;Љl$������l$��u<���   �@�FD�����   �D$P�@�FD�\��VH���   �:���   @���   ��u{���d$(����!����t%�D$P�d$,����!����t�VH�:�:�P�A���   �VD�D$(�@�����   �VD�D$,�@�\��FH���   �T8���   @���   ����   ���d$4����!����t#�D$P�d$8����!����t�FHǋ�P�|�D$(�d$4����!����t$�D$,�d$8����!����t�FHǋP�P�A���   �VD�D$4�@�����   �VD�D$8�@�\��FH���   �T8���   @���   ���  ���
  �d$@����!����t&�D$P�d$D����!����t�FHǋ�H��   �D$(�d$@����!����t)�D$,�d$D����!����t�VH�L:�:�H�   �D$4�d$@����!����t&�D$8�d$D����!����t�VH�L:�:�H�V���   �D$@�@�FD�����   �VD�D$D�@�\��FH���   �L8���   @���   ��VH�؋L:�:�H��؋FE��;�l$��������   3�;É\$��   ���  �nd�VD�����D��\$� �$h8W�3�  ����W��S  ���   B���   �?u=���  t4���   �D$ 3��L$�D$$�D$�l$ �t$��!��  P��{  ���D$���   @��;��D$�g������   ���  Rh�7W覔  ���NdW�ZS  �D$P�h  ���   ][_^��x� ����������������DSUV��W�~���;�v���T$X3ۉ^0�lyShO  �HHR�Qx��;�u_^]3�[��D� ���te  ��ly�S�HS��R��H  ��;ÉF,uh�8�w`  ��3�_^][��D� �ly�VSS�H��R��H  ��;ÉF0uh�8�=`  ��3�_^][��D� �F�\$X;���  3ɋ��  ���E �*  �U���D$�D$�E��!�T$���D$�D$����!�\$L�D$�U ��!�E���\$P�T$���D$�U��!�\$$�D$���D$�T$����!�\$(�D$�E ��!�U���\$,�D$���D$�E��!�\$0�T$���D$�D$����!�\$4�D$�U ��!�E���\$8�T$���D$�U��!�\$<�D$���D$�T$��!�\$@�D$��!���-  �U�D$���D$�T$����!�E ���D$�U��!�D$�������\$L�D$�T$�E ��!�\$P�D$�D$����!�U ���\$$�D$�E��!�T$�������\$(�D$�D$�U ��!�\$,�D$�T$����!�E ���\$0�D$�U��!�D$�������\$4�D$�T$�E ��!�\$8�D$�D$��!���\$<�D$��!���U�\$@���T$�D$��!�F$����l$�\$D�X�P�F+����3���3҃�;���  �É|$���D$�n,�D$���uV�E ������!����tB�E�d$L����!����t,�E�d$P����!����t�F0���<���   H���   ��uY�E �d$$����!����tC�E�d$(����!����t-�E�d$,����!����t�F0���|���   H���   ��uY�E �d$0����!����tC�E�d$4����!����t-�E�d$8����!����t�F0���|���   H���   �D$��t^��uY�E �d$<����!����tC�E�d$@����!����t-�E�d$D����!����t�F0���|���   H���   ��+�t�l$�FG��;��l$�]����l$��u>�F�~,�@���F�~,�D$L�@�\��F�~,�D$P�@�\��F0�~�<�F@�F����   ���d$$����!����t:�D$L�d$(����!����t#�D$P�d$,����!����t�F0��8�x�C�F�~,�D$$�@���F�~,�D$(�@�\��F�~,�D$,�@�\��F0�~�|�F@�F����   ���d$0����!����t=�D$L�d$4����!����t&�D$P�d$8����!����t�F0��8�x�   �D$$�d$0����!����t;�D$(�d$4����!����t$�D$,�d$8����!����t�F0��x�x�C�F�~,�D$0�@���F�~,�D$4�@�\��F�~,�D$8�@�\��F0�~�|�F@�F���G  ���M  �d$<����!����t?�D$L�d$@����!����t(�D$P�d$D����!����t�V0�
�
�P��   �D$$�d$<����!����t>�D$(�d$@����!����t'�D$,�d$D����!����t�F0��P�P�   �D$0�d$<����!����t;�D$4�d$@����!����t$�D$8�d$D����!����t�F0��P�P�V�F�V,�D$<�@���F�V,�D$@�@�\��F�V,�D$D�@�\��F0�V�T�F@�F��F0��؋P�P��؋D$X�V@��;D$X�l����F�D$X    ����   ���  �^d3�F,��Ń����@�\$�@�\$� �$hh8W迋  �� ��W�tJ  ���   B���   �?u=���  t4���   �D$3��L$�D$ �D$�l$�t$��!衍  P�gr  ���D$X�N@��;��D$X�b����V���  RhP8W�8�  ���NdW��I  _^]�   [��D� �������������U������L  �lySV�uW3���W�HHh�  V�Q|�ly�D$ h�  V�BH���   ���L$0�D$��n  �ly�|$Wh�  �QHV�|$(�R|�C$�lyh�  V�HH���   �C�ly���΋��   �PxP�L$4�\o  ���  jh   V�L$<�ep  �����3����I�����|$~�d���+ˊ< t<	u�_F�1;�|�D$0�L$HPh`9�n  �L$$PQ�Uo  P�q  ���L$ �n  �L$H�n  �u<��tQ��  ��tG�����3��ly�D$�R��Ij j �LQ��H  �����  �D$QVhX9P藉  ���A�lyj Gj �BW��H  �Ѝ��  ���3����T$���+����������ȃ�󤋃�  ��t;��  ��t1��  ��t'�sdhT9����G  �L$Q����G  hP4����G  ���  ��t=��  ��t3��  ��u)�sdhL9���G  ���  ��P�G  hP4���G  �D$���  �T$�D$�z�E0�O�E�O����  �D$D    �D$@�����E$������  �����E�E4�O�E�O����E(����E�E8�O�E �O����E,����E�l$X�\$,�t$,���\$�t$,�\$�t$,�$h49V��  �� �KdV��F  ���   B���   �?u=���  t4���   �D$H3��L$ �D$L�D$$�l$H�t$ ��!���  P��n  ���D$��H�D$������D$P���  h 9V蕇  ���{d��V�GF  ����E  �T$3���lyWW�H�C����R��H  �s4��;ǉu+h9��S  �D$P�g  ���L$0��k  3�_^[��]�8 ���  h 9$�L$$���  �{�{�{�k  P�n  ���L$ �k  �L$�UQR����G����uA�D$P�Bg  ������������������*���V�$g  ���L$0�>�fk  3�_^[��]�8 �C���   ;�t9��  t�u��V������u���   ��u�C�{;�t9��  tV���������u�{9{uI9��  t<�L$�T$QR�D$`h�8P�%�  ���L$XQ�L$$�j  P��e  ���L$ ��j  9{t9��  t�T$��RV�����D$�D$���   ���   �S���   ȉ��   ���   �D$��P���   ���   �f  ���������L$0�Pj  �D$_^[��]�8 ������   SUV3�W��Vh  �?V��$�   �l$`�K  h  �?VV��$�   �8  ��$�   �|i  ��$�   �t$�t$��R  ��$  ;���  �ly��$�   SR�HH�Q@�   ���|$$���3��L$XW��  �D$$،$0  �D$ ،$$  ��ل$  �L$��؄$  �\$Xل$4  �L$$ل$(  �L$ ��ل$  �L$��؄$  �\$\ل$8  �L$$ل$,  �L$ ��ل$   �L$��؄$  �\$`�D$0،$0  �D$,،$$  ���D$(،$  ���\$d�D$0،$4  �D$,،$(  ���D$(،$  ���\$h�D$0،$8  �D$,،$,  ���D$(،$   ���\$l�D$<،$0  �D$8،$$  ���D$4،$  ���\$p�D$<،$4  �D$8،$(  �lyWh�� S���D$@،$(  �HH�|$X�|$\��ٜ$�   �D$H،$D  �D$D،$8  ���D$@،$,  ��ٜ$�   �D$T،$<  �D$P،$0  ���D$L،$$  ��ٜ$�   �D$T،$@  �D$P،$4  ���D$L،$(  ��ٜ$�   �D$T،$D  �D$P،$8  ���D$L،$,  ��ٜ$�   �Qx����;���   ��$�   �fP  �ly��$�   QV�B@�P`����$�   ��$�   R�zP  ��$�   �P  ��$�   ��$�   P�P  ��$�   �P  Wh�  ��$�   �Q  ;ǉD$LtWh�  ��$�   ��P  �D$P���T  �ly���|$���   ���R=�  ��   ��$D  ��t5���  �ly���   �Rxj���  h   Q����g  ǅ�     �@�6���3�ǅ�      ���+����  ���������ȃ��|$ǅ�      �D$L��u@��t��u7��$<  ��t,��$@  �t$XQ�   ��0���S���)�������  �|$��$<  ���I  �   �F  �ly�ˋ��   �P=  uϋly���   ���RxP��$�   ��e  ���  jh   V��$�   ��f  �����3����I�х�~�d�����+̀8 u� _@�<;�|���$@  �ly��t@�h���3�j ���Ij �LQ��H  ��$L  ���D$VRhX9P�R�  �l$d���7�Hj Bj R��H  �Ћ����3����T$���+����������ȃ�󤋌$D  3��L$�ly��Ph�  �JHSF�Qx���������j ���KQ  �D$�Ѓ�u3��D$P��u7�ly�ˋ��   �P4�L$�T$QRV�   ��0��$�   ���P�������ly�ˋ��   �R(�؍D$3�P�t$��_  ��;މt$�E�����D$��t�L$Q�_  ����$�   �D$    �sM  ��$�   ��c  _^][���   �@ �����������T$���L$��L$�P�H� ���������� �������������DSUVW�ك��̉\$,���  �kdP�oj  ���<  ����  h�9�L$�2c  P�e  ���L$�Pc  ���  �n  P���7���H3���3��Ü  ���+�S�ы������ʃ����=  ��2���3�S���+����������ȃ�����<  ��9���3�S���+��ы������ʃ����<  �p9���3�S���+����������ȃ����<  ��2���3�S���+��ы������ʃ����e<  ��2���3�S���+����������ȃ����;<  ��2���3�S���+��ы������ʃ����<  ��2���3�S���+����������ȃ�����;  �H3���3����+��ы������ʃ�S���;  �\$���  ��t���hf���D$    �L$�D$    �D$�D$    �T$�L$(�D$    �L$�D$$�T$,�D$  �?�D$�D$    �T$�L$4�D$  �?�L$j �D$4�T$<�D$    �D$�D$     �T$ j �L$H�D$     �L$ j�D$H�T$P�D$     �D$ �D$(  �?�T$(��0��$�   �   �t$`����$�   ��$�   󥋋�  �l  P���v������:  �Kt�w:  �KP��@  _^][��DÐ��������H  �L$ ������$L  j �Sm  ����$�  ��   j���k  P�L$(�2����tph:�L$�`  �D$ ��$�  Pjj�Zg  ��t@h:�L$��_  P��$�  ��h  �L$�`  �L$ Ǆ$�     Q��-������u�L$ ��_  �L$ �$���3���H  � j�Ba  ����a  �L$ ������a  j�%a  ���L$ �_  �L$ ������   ��H  � ���   @� ���������� Vj�ur  ���L$P��^  �L$��_  ��u�L$�B_  �   ^�� �j j j�m[  ������t���-p  ��!�3�h�p�L$��^  �D$VP����h :��^  �L$j Qh�� �m  ��$�L$����^  �L$��^  ��^�� ÐÐ��������������SUV��W�~t���P;  ���   ���C;  ���   �8;  ���   �-;  ���   �";  ���   �4  ��  ��d  3ۋω�^�^�^�^�^�^�^�^ �)@  ���"@  ���   �W>  ���   �L>  ���   �A>  ���   ���   ���   ��   ��  �^�   ��,  ��8  ��<  ��@  ��D  ��H  ��L  ��P  ��T  ��X  ��\  ��`  ��t  ��x  ��h  ��l  ��p  ��|  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ǆ0     ǆ4  �  �^H�^L�^`�^d�^P�^T�^\�^X�^h�^l�^p��  ��_^][Ð����������������SUV��NHW�FH��t	P�wX  ���NL�FL��t	P�dX  ���N`�F`��t	P�QX  ���Nd�Fd��t	P�>X  ���NP�FP��t	P�+X  ���Nl�Fl��t	P�X  ���Nh�Fh��t	P�X  ���Nt�L$ �6>  ���   �L$�'>  ���   �L$�X<  ���   �L$�I<  ���   �L$�:<  �Np�Fp��t	P�W  ���FT�nT��t5�N3ۅ�v#�x�G���t�? t	W�W  ���F��C;�r�U�kW  ���FX�nX��t5�N3ۅ�v#�x�G���t�? t	W�@W  ���F��C;�r�U�,W  ���F\�n\��t;�N3ۅ�v)��x  �G���t�? t	W��V  ���F�ǀ  C;�r�U��V  ����  �Ib  ���   �1  �L$��7  �L$��7  �L$��7  �L$�z;  �L$ �q;  _^][��Ð����������  �vx  U��3�h   ���   h�p�D$���   �2  ���,  S�\$VW���   �D$,    B�D$(    ���   �D$$    ��p��݃�S�  3Ɋ���$�`�=�p ��   �=�pr��   �=�p ��   �T$TRh`;h�p�u  ������   h�p�A  �����3������+��T$T���������ȃ�󤋍,  ��@��,  �L$TQ���   �6  �E�]��  ShT;h�p�=u  ����u;h�p��@  �����3������+��ы������ʃ�󤋅,  ����,  �\$h   h�p���   �?1  �������_^��[��  �}  ��  �   ]�Ĵ  � ��p< ��   <nt@<tu��D$(�L$$PQhH;h�p�t  ����u���,  �E��@��,  �E�n����T$,�D$(R�L$(PQh<;h�p�Ft  �����D�����,  �E��@��,  �E�)����T$,�D$(R�L$(PQh0;h�p�t  �����������,  �E ��@��,  �E �������$T  Rh(;h�p��s  ���������h�p�?  �����3������+���$T  ���������ȃ�󤋍,  �� ��,  ��$T  Q���   �4  �E�d�����$T  Rh;h�p�Cs  �����A�����,  h�p�π   ��,  �?  �����   P�Z4  �E�����D$PPh;h�p��r  ���������p��p<ot��p�E��uh;���   �4  �E�E��uh�:���   ��3  �E�E��uh6���   ��3  �E�L$H�T$Q�D$HR�L$ P�T$LQ�D$$RPh�:V�^r  �� ��u`��u	�   �\$h�4V3��xs  �����  ��$T  �NQVh�:P�r  ����uG��h�4j �>s  ����u��  �T$H�D$8R�L$ P�T$LQ�D$@R�L$(P�T$TQ�D$HR�L$0PQh�:V�q  ��,��	ud��u	�   �\$h�4V3���r  �����y  ��$X  �V�N�RVQh�:P�vq  ����uG��h�4j �r  ����u��  �T$8�D$R�L$8P�T$ Q�D$<R�L$$PQh�:V�)q  �� ��u`��u	�   �\$h�4V3��Cr  ������  ��$T  �VRVh|:P��p  ����uG��h�4j �	r  ����u��  �D$�L$P�T$QRhl:V�p  ����u\��u	�   �\$h�4V3���q  �����b  ��$T  Vhh:P�gp  ����uG��h�4j �q  ����u��
  �D$�L$P�T$QRhT:V�)p  ����u\��u	�   �\$h�4V3��Cq  ������   ��$T  Vhh:P��o  ����uG��h�4j �q  ����u��   �D$8�L$P�T$8Q�D$ R�L$<P�T$$QRh8:V�o  �� ���������u	�    �\$h�4V3��p  ����tW��$T  �NQVh,:P�Xo  ����uG��h�4j �|p  ����uу�vWW�Mt�84  ��t�E �E���ǉE�E����3�]�Ĵ  � ��t� z �� � ^  �� l�  ��������������SUV��W�F��tJ��,  ����j ��,  �ly���Qj P��H  ���FP��uh9�c:  ��3�_^][��ËF ��t[3�3ۅ�v3S�Nt�^4  ����t�O�WQR���   �3  �;�v��F C;�r͡lyj ��    j �HR��H  ���Fp�F��u�F   �F��t;�ly�@j j �Q��P��H  ���F`��uh�;�9  ��3�_^][��ËF��t;�ly�@j j �Q��P��H  ���FL��uh�;�o9  ��3�_^][��Ë��t;�ly�@j j �Q��P��H  ���FH��uh�;�.9  ��3�_^][��ËF����   �lyj j �Q��    +���Q��H  ���FT��uh�;��8  ��3�_^][��Ë��F3ۅ�vA���   j jW��L  ����S��0  P�L$�P  P���Q  �L$��P  �F��C;�rŋF����   �lyj j �J��    +���R��H  ���FX��uhx;�J8  ��3�_^][��Ë��F3ۅ�vA���   j jW�BL  ����S�G0  P�L$�P  P���uP  �L$�<P  �F��C;�rŋF���  �lyj j �Q�@����P��H  ���F\��uhh;�7  ��3�_^][��Ë؋F3���vQ��`  j h�  S�K  �����   W�/  P�L$�O  P����O  �L$�O  �F�À  �ŀ  G;�r��ly�Fj j �Q��P��H  ���Fh��u_^][��Ëly�Fj j �Q��P��H  ���Fl��u_^][��ËNj ��QP�K  ��_^]�   [��Ð������SVWj j �>  ���D$���8  �}K  ���D$�  �L$j Q����K  ����   �\$�lyj j �B��    Q��H  ��3��ۉD$~,�|$ �T$�L$WR�L  �L$���D$�<� tOF��;�|؋T$�L$j SPR�L  ���D$P�J  ����uN�L$Q�=  �T$R�
K  ��3�_^[��� �T$R��I  �D$P�x=  �L$Q��J  ��3�_^[��� �L$j j j �1K  ��t�t$�T$R�J  ����_^[��� �D$P�'=  �L$Q�J  ��_^3�[��� �����������������S�\$UV��W����  �ly�[j j �H��R��H  ���D$$����  ��v=�T$(3��\$�
�nHǃ��I���L� �)�(�i�h�I�H�D$H�D$�D$$u�PS���������D$u�T$$R�H  ��_^][���  �lyj h�  P�QH�R|�T$(��lyh�  R�HH���   �����F@�NtP�.  ���D$tH3ɉx��v?�T$(�T���T$��\  �@��t	�T$(����T$����T$�D$A��;ˉT$rͅ���  �L$4�߃� �����D$    �T$4�l+��|$�l$��\  ��u�Ջz�j3�;��*�Ã����\$(���,��i��j�,��)�j�,��iu�j��j��3�Y�\$,;�t9�*���,��i�j�,��i�j�,��iu�j��3�Y��j��3�Y��i�i�i�i�\$0;�t9�*���,��i�j�,��i �j�,��i$u�R3���Q(��R3���Q(��i�i �i$�i(�T$<�ZC�Z�T$8�ZC�Z�T$@��p  C;ŉ�p  �V,�Q��V(�Q�V$�Q�V<�Q�y,t%�x�T$�^<����T$�V,�P�V(�P�V$��~<�T$4�l$G�~<�|$��P����O�T$4�l$�|$�|����^@�D$CP�^@�:  �L$(Q�MF  ��_^][���  �L$(�D$4����P�Q�P �Q�P$u�I��I�H(�L$,3�;�t&�9���x,�y�x0�y�x4u�I�H8��I�H8��P,�P0�P4�P8�L$0;�t&����P<�Q�P@�Q�PDu�I�HH��I�HH��P<�P@�PD�PH�L$<�iE�i�L$8�yG�y�L$@��p  B��p  �N,�H�V(�P�N$�H�V<�P�XL�F<_^][���  ��� 2  �6g  U��3�h   �MT�UX�L$�M\�L$���   h�p�E0�E4�E8�E<�E@�E$�E(�E,�T$���   �9!  ����	  SVW���   B���   �?u4���   �D$ 3��T$(�D$$�D$,�l$ �t$(��!�tf  P�:K  ����p��݃�S�f	  3Ɋ���$���=�p �J	  �=�pr�=	  �=�p �0	  �T$0Rh`;h�p�,d  �����	  h�p�0  �����3������+��T$0���������ȃ��L$0Q���   ��'  ��    �E,+ЋEX���L$�  ��p< �  <n��   <t��  �E8�M;���  �@�E`���HQPhH;h�p�}c  �����a  ��t  ��t�E8�� �@�E`�$������x  ��u�E8�U`�� �@�d��D���E8�M`�@�D�  �?�E8@�E8�   �E4�M;���  �@�EL�4��~�^WSVh<;h�p��b  ������  ������\  ��t������������E4�  �E4@�؉E4�  �E0�M ;���  �UH�@�4��~�^WSVh0;h�p�pb  �����T  ۅ4  ��ۅ4  ����4  �؉D$�D$���E0�$  ��$0  Qh(;h�p�b  �����  h�p�e-  �����3������+���$0  ���������ȃ�󤍌$0  Q���   �%  ��    �E(+ЋET���L$�  ��$1  Rh;h�p�a  �����}  h�p�-  �����   P�b%  �@�E$���M\����D$�J  �E<�M;��<  �MP����پ�p�    ��p<ot��p��$ 
  ��$
  R��$
  P��$
  Q��$
  R��$
  P��$
  Q��$
  R��$
  PQh�:V��`  ��,��	��   �h�4���V3����a  ����t:��$
  �V�N�RVQh�:P�`  ����uG��h�4j �a  ����u�3Ʌ�vJ��$
  �B���}E0�H���0  ���}E8�H���p!  �B��}E4�H���@)  A��;�r��T$�D$�L$RPQ��$L)  S��$�!  RP��  ��$
  ��$
  R��$
  P��$
  Q��$
  R��$
  PQh�:V��_  �� ����   �h�4��@V3����`  ����t6��$ 
  �VRVh�:P�_  ����uG��h�4j �`  ����u�3Ʌ�v6��$
  �B���}E0�H���0  ���}E4�H���@)  A��;�rыD$�L$�T$PQR��$L)  SP��  ��$
  ��$
  R��$
  P��$
  Q��$
  R��$
  PQh�:V��^  �� ����   �h�4�ʀV3����_  ����t6��$ 
  �VRVh|:P�^  ����uG��h�4j �_  ����u�3Ʌ��  ��$
  �B���}E0�H���0  ���}E8�H���p!  A��;�r���   ��$
  ��$
  R��$
  P��$
  Q��$
  R��$
  PQh8:V��]  �� ����   �h�4�ʀV3���_  ����t6��$ 
  �VRVh,:P�]  ����uG��h�4j ��^  ����u�3Ʌ�v6��$
  �B���}E0�H���0  ���}E8�H���p!  A��;�rыD$�L$�T$PQRS��$�!  j P�  ��$
  ��$
  R��$
  PQhT:V�]  ������   h�4V3��>^  ����t2��$ 
  Vh�;P��\  ����uG��h�4j �^  ����u�3Ʌ�v��� 
  ��}E0�H���0  A;�r�T$�D$�L$RPQSj ��$D  j R�m  ��$
  ��$
  P��$
  QRh�;V�b\  ������   h�4V3��]  ����t2��$ 
  Vh�;P�/\  ����uG��h�4j �S]  ����u�3Ʌ�v��� 
  ��}E0�H���0  A;�r�D$�L$�T$PQRSj ��$D  j P�   ��$
  ��$
  Q��$
  RPhl:V�[  ������   h�4V3���\  ����t2��$ 
  Vhh:P�v[  ����uG��h�4j �\  ����u�3Ʌ�v��� 
  ��}E0�H���0  A;�r�L$�T$�D$QRPSj j ��$H  QW�������h   h�p���   �Y  ���#���_^[�U@�E<�U �E�   ]�� 2  Ð�.��R ����������SUVW����̍�  ���   P�E  ���)  ��3�;�th8<��&  ����_^][��� ���   �  ���   �  ���   �  h$<�L$�)>  P�@  ���L$�G>  �L$$Q���[�����uh<�&  �������_^][��� h <�L$��=  P�g@  ���L$��=  ��������u�����_^][��� h�;�L$�=  P�-@  ���L$��=  ����  ����������u!��  h�;�^%  �������_^][��� ��  �N�FT3�;�v:�x9/t%�ly�UU�B��Q��H  ��;ŉG�D  �o�F��C;�rɋN�FX3�;�v:�x9/t%�ly�UU�B��Q��H  ��;ŉG��   �o�F��C;�rɋN�F\3�;�v@��p  9/t%�ly�UU�B��Q��H  ��;ŉG��   �o�F�ǀ  C;�rƋV�FP3�;���   �P�B���P�<�    +��FT�\����x���hE�h�B��<�    +��FX�\����x���hE�h�B��<@���~\��ǋ�t  ��x  ����t  EA��t  �F;�r����WI��3�_^][��� h�;��#  �������_^][��� �����������������T  �D$TSVW��jh   �L$��  PQ���GD  ��� =  �L$�;  �|$`���3��T$`���I����D$`P��������t.hH<�L$�A;  P�6  ���L$�_;  _^3�[��T  � ��8  ����   �F  ������   �L$(��A  �L$D��A  �L$Q����B  P�L$H�,D  �L$�#B  �T$��R�'C  P�L$,�D  �L$�B  hD<�L$�:  P�L$,�C  �L$��:  �D$(��P��F  �L$DQ���G  W�UG  ���L$D�A  �L$(�A  ���$d  ��@  ��t�T$`��RW� o��_^�   [��T  � ��D  ��t�D$`��PW�h}��_^�   [��T  � ��H  ��t�L$`QW���Ћ��_^�   [��T  � �T$`��RW��f��_^�   [��T  � ����  �L$ V�0���h�<�L$�9  �D$��$4  Pj j��@  ����   h�<�L$�w9  �L$Q��$8  �vB  �L$���9  ��tRj� ;  ��$�  ���L$$R�<D���;  j ��;  j��:  ���L$�M9  �L$$�d����   ^���  � Sh�<�L$��8  �D$��$8  P��A  ���L$���9  ��[t"hT<�L$��8  P�4  ���L$��8  ��L$$Q�:������u�L$��8  �L$$�����3�^���  � j�*:  ��$�  ���L$$R����j ���;  �:  j�:  ���L$�u8  �L$$������^���  � �� Vj�eK  ���L$P��7  �L$�8  ��u�L$�28  �   ^�� �j j j�]4  ������t���I  ��!�3�h�p�L$��7  �D$VP����h�<�7  �L$j Qh�� �F  ��$�L$����7  �L$�7  ��^�� ÐV����H  �D$t	V�4  ����^� ��SVW���.  �~���,  �^,���"  �N@�K  �NL�K  �L$�D$�N`����!�FX�w  ���p  �+=  �F\��_^[� V���   �D$t	V�3  ����^� ��SV��W�~��!���+  �^,���!  �F\P��<  ���NL�mK  �N@�eK  ���  ���  ���-  _^[Ð�����������VW����,  �F`j j P���x,  ����tj-V�N@�J  j.V�NL�|J  ��_^Ð��������V��F\��tOP�N@�D$+   �D$    �K  P�D$P����)  �N\�D$,   Q�NL�D$    �K  �T$PR����)  ^��Ð����������������  SV��L$4��  �L$H��  �L$��  �B  ��t/���A  �؅�t"�ly�ˋ��   �R=�  u����+  ��u&�L$�  �L$H�  �L$4�  ^3�[�Ĕ  �UWhtxt heman�L$�X!  �D$�N@Pj��I  �L$(�P  P�L$��  �L$(�  htxt heman�L$�!  �T$�NLRj�I  �L$(�  P�L$@�  �L$(�  �L$(��  P�L$T�|  �L$(�c  ��$�   �W4  �L$t�N4  3��ly��Ph)  �QHSG�Rx����tK�ly���   ���RxP��$�   ��4  j��$�   h�   P��$�   ��5  ��$�   Q�N�F  똋NXj h�  �  3�3����D$��   �^�L$d�3  �NXP���  ��$�   RP�a  P�L$x�G4  ��$�   �4  �L$d�4  j��$�   h�   Q��$�   �75  ��$�   ��R��  ���t!��$�   �N,P�  ��$�   ��Q���2  �D$G;��c���3�����   W�N,���  �|  P�L$h�R3  �NXPS��  �L$d�o3  �L$(��2  �NXP��$�   SR�  Pheman�L$X�  ��$�   �93  �L$(�03  �D$P�NLPW��G  G;�|��D$;�}�����  Q�NX��  �D$G;�|�NXUh�  ��  �^���  ��3���~=W����  P�L$,�2  Pheman�L$D�
  �L$(�2  �T$<�N@RW�sG  G;�|Í~@���4F  �^L���*F  jj����G  jj����G  ��������L$t�d2  ��$�   �X2  �L$��  �L$P��  �L$<�  _]^�   [�Ĕ  Ð�������������D$��  HSUV��-W����  3Ɋ��)�$��)�F\���n  �^@P���AG  ���[  �L$�P1  �L$,��  �N,�o  �N\��T$�D$RPj �D$     ��7  ����   �D$�L$;���   �~�L$,QP���yF  �L$@��0  P�T$themanR�L$8�  P�L$ �1  �L$p�I1  �L$@�@1  j��$�   h�   P�L$(�x2  ��$�   Q���)  ���t<�T$��R�8F  ��$�   ��P�y  �L$,��QP�NLE�E  ��$�   �N,R�  �D$�L$@;��D$�=����D$�L$�T$@Q�N\RP�D$ ��6  ���������8D  �NL�0D  �L$,�  �L$�~0  ������_^]�   [�Ā  � �F\���t  �^LP���E  ���a  �L$�/  �L$,�5  �N��
  ��D$�L$PQ�N\j �D$     �O6  ���   �D$�L$;���   �~,�T$,��RP��D  ��$�   �[/  P�D$dhemanP�L$8�  P�L$ ��/  �L$`�/  ��$�   �/  j��$�   h�   Q�L$(��0  ��$�   ��R�  ���t<�D$��P�D  ��$�   Q����  �T$,��RP�N@E� D  ��$�   �NP�   �D$�L$@;��D$�7����D$�L$�T$@Q�N\RP�D$ �O5  ��� ����N@�B  ���B  �L$,�o  �L$��.  ���o���_^]�   [�Ā  � �NXj h�  �  �n,�D$���`	  ��3���~0W���  P�L$T�f.  �NXP���  P��  �L$P�}.  G;�|Ћl$;�}�����  Q�NX�/  G;�|�NXSh�  �<  _^]�   [�Ā  � ��)�%k'�(�) ��������dS�\$pV�t$pW����u_��t[�lyV�H@�Qh����tHj)P�L$�(���j j j�j��L$�w$  ���L$u����_^3�[��d� �z���_^�   [��d� �T$|��RSV�C  _^[��d� �������0j�f@  ���L$ P��,  �L$ ��-  ��u�L$ �3-  �   ��0�Vh�<�L$(��,  h�p�L$��,  �D$$j �L$PQh+�T$jRh�� �+D  ���L$����,  �L$$��,  �L$��,  ��^��0Ð���Vj j j��(  ������t���=  �"��^�3�^Ð������ly�T$R�H@�Qh����j h�  �?  �   � ���������dS�\$pV�t$pW����u_��t[�lyV�H@�Qh����tHj*P�L$����j j j�j��L$��"  ���L$u�����_^3�[��d� �����_^�   [��d� �T$|��RSV�A  _^[��d� �������0j��>  ���L$ P�Y+  �L$ �0,  ��u�L$ �+  �   ��0�Vh�<�L$(�[+  h�p�L$�M+  �D$$j �L$PQh�,�T$jRh�� �B  ���L$���M+  �L$$�D+  �L$�;+  ��^��0Ð���Vj j j�d'  ������t���$<  �X"��^�3�^Ð������ly�T$VR�H@�Qh������jh�  �  jh�  ���  �   ^� ������lyVW�|$��W�H@�Qh�T$�D$����RPW�G@  _^� ����0j!�=  ���L$ P�*  �L$ ��*  ��u�L$ �c*  �   ��0�Vh =�L$(�*  h�<�L$�*  �D$$j �L$PQh�-�T$jRh�� �[A  ���L$���*  �L$$�*  �L$��)  ��^��0Ð���Vj j j�$&  ������t����:  ��"��^�3�^Ð�����V��3���F�F�F�F�F�e3  �F��^Ð���������������Q�W3  YÐ����V��F�F    ���F   t �lyj j h   �H��H  �����u�L$�_0  �����^� �Nh1D4ChCD4Cjj �T$jR�	3  �N��u�3  �L$���"0  ��^� �3  �L$�F�F    �0  3�^� ��������������V��j j �N�A3  �F   �F    ^ÐV��N��2  �> t	V�J$  ���    �F    �F   �F    �F    ^Ð��V��W�N�F;�|_3�^�+�=   }�F��F   �~���j PQ�N�e2  ;�}�F   _3�^ËF�F    �_�F�^ÐQSUV3�2�W�|$��\$�\$�E�M;�|���x�������   �M�U �A<
�MtK<tG<\u�L$��u�D$�D$뺄�u< t�<	t���u	<#u�D$�>�D$FH;��D$ t=닊D$�D$ ��t&���v����|>� �k����L$�> FI;�t�X������P����> ��_^][Y� �����������V���F    �F    ��0  �F�lyj j �Hh  ��H  �����^Ð������V��F��t�   �N�F    ��t�> u�L$��-  �����^� h1D4ChCD4Cjj �D$jP�0  ��u�N�F1  �L$���-  ��^� �L$�F   �-  3�^� ���������������V��W3��N;�t9~t�F;�t	P�P�0  �~_^Ð�������V��F��t�F��t�����N�20  �F    ^Ð��������V��W�|$�> t*�? t%�F����F@G=   �F|���n����? u�_^� ����V��F��t�����> t	V�V!  ���    ��V�d/  ���    ^Ð���������T$���L$��@    �P� ��������;   ������������Ð�������������AÐ������������AÐ������������3�;�Vt�q�p�A;�t�1�0��Q^Ð��������������V��Wj �~j ���^����    �~�    �F    �F    ��_^Ð�����������V���   �N�@���^Ð��������������AÐ�����������V��j�   ����t"�L$�VQR��������N�A�A�F�^� �N3��A�A�F�^� ���������V��W�|$;~u
��������F�F;�t���tH���t������W�h   ��_^� SV���W�������t.UW�k������;���t��t���d���V�.   ������u�_]�C�    �C    �C^�     [Ð������VW3��W�����t�|$;�s���4���F��u�_3�^� ��t����-���_^� ��������V���X�����^Ð���V���h  ������^Ð��������������SUVW��������l$����tG���������t/�����:u��t�P��:Vu������u�3��������tW����������u��ly�����j �P3����j Q��H  �Ћ����3������+�R���������ȃ�����������#���_^][� ������������QSUVW���D$ �����l$����tG��������t/�����:u��t�P��:Vu������u�3��������th�����������u��ly�����j �P3����j Q��H  �Ћ����3������+�R���������ȃ����4����D$_^]%�   [Y� �D$_�D$^]%�   [Y� �������������QSUVW���D�������tl�l$���3������D$t/�����:u��t�P��:Vu������u�3��������t�����������u�_^][Y� �D$P�  ����W�����_^][Y� ����������SUVW3���������tL�\$��������t/����:u��t�P��:Vu������u�3��������t��E�Y�������u�_^]���[� _��^][� SUVW3��E�������tL�\$���4�����t/����:u��t�P��:Vu������u�3��������t��E���������u�_^]3�[� _��^][� �VW3��������t�|$;�t��F������u�_3�^� ������_^� ������������QVW����������t)���������D$t�D$P�W  �����]�������u׋�����_^YÐ�����������V���h  �������^Ð��������������Q�lySVW��j �Hj j ��H  ���D$��tA�|$�lyj j �B�4�    V��H  �L$���A�D$�H��u�T$R�  ��_^3�[Y� �x�lyj j �HV��H  �T$���B�D$�H��u��P�m  �D$P�c  ��3�_^[Y� �t$�lyj j �Q��    P��H  �L$���A�D$�H��u,��P�  �T$��R�  �D$P�  ��3�_^[Y� �p�L$Q�������D$_^[Y� ��������������D$P����� ���QVW�����������tj����������D$tN�P�H��tQ�  �D$���P�H��tQ�z  �D$���H����t	P�c  ���D$P�V  �����\�������u�������_^YÐ������������   V��F����   ��$�   SP�L$�*  P�L$,�$  h=�L$�  P�L$H��#  �vj �L$,j��T$LQ��$�   RP��'  ����$�   PQ�I&  ���T$lPR�;&  ����P�p  ���L$`���$  �L$|��#  ��$�   ��#  �L$D��#  �L$�  �L$(��#  �L$�  ��[u�   ^�Ĭ   � 3�^�Ĭ   � ��������V��F��tR�lyWP�Q�R�ly���F�QP�R�L$ ���T$h  WP�D$j +�j Q�L$$+�RP�FQP���  _^� �ly����yV�0��-  ��u^��Á�@  }3�^����~�����u^���������u^���������u^����4�����u^����V�����u^���h�=�L$�o  �L$Q�  ���L$�  h`=�L$�K  �T$R�a  ���L$�e  h=�L$�'  �D$P�=  ���L$�A  h`=�L$�  �L$Q�  ���L$�  h�=�L$��  �T$R��  ���L$��  �   ^��Ð�����������������������������������������h�   h�xh�� �l  ����tk��xHtHHtHu<��x   ���x   �   �dy�hyh�   h�xh�� �N  ����xø   ��x   �\y�`y�VW��=���3���x   ���+�h�   ������xh�x���ȸ   ��h�� �3���x�  ��x��x��x� y�y�y�y�y�y�y�y�$y�(y�,y� y�0y�4y�8y�<y�@y�Dy�Hy�Ly�Py�Ty�Xy�\y�`y�dy�hy�3  ����x_^Ð�������h�   h�xh�� �  ��Ð��������D$����tE�8 t@�QA��u�I;�t�9 t���	t
��
t��u� �����t�� t��	u�H@��u�ËD$P��������t1���t+VW�   3���+���:t
��/t��\u�<�JB��u��_^Ð�������������D$P�V�������t�8 t�Ȋ�� t��	u�_�QA��u�Ã�0�L$ V�t$8V��  Ph�=�L$��  P�D$P�  P��  ���L$�  �L$��  �L$$��  V�L$�  Ph�=�L$�  �L$(PQ�\  P��  ���L$$�  �L$�  �L$�  ^��0Ð����0�L$ V�t$8V�^  Ph>�L$�O  P�D$P�  P�^  ���L$�b  �L$�Y  �L$$�P  V�L$�  Ph >�L$�  �L$(PQ�  P�F  ���L$$�  �L$�  �L$�  ^��0Ð���lyV��Hj�V���   ����^Ð�����T$�lyV��HRV���   ����^� �lyV��Hj�V���   �ly�L$�Bj VQ���   ����^� �������������ly�PQ�RYÐ��ly�T$V��Hj VR���   ����^� ���������������ly�PQ�R��ály�P�D$PQ�Rh��� ����������ly�P�D$PQ�Rl��� ���������VW�|$��W��������u	�D$_^� �ly�HWV�QH��_^� ���������������VW�|$��W�������u	�D$_^� �ly�HWV�QL��_^� ���������������VW�|$��W�R������u	�D$_^� �ly�HWV�QD��_^� �����������������VW�|$��W�������u"�L$ �1�D$�Љ2�q�r�I_�J^��� �ly�BW�L$VQ�P`�Ћ2�D$$�ȉ1�r���q�R_�Q^��� ����VW�|$ ��W�������u�D$$�t$P���:  _��^��� �ly�QWV�RP���L$�D$ ��  �D$ ��t
P�L$�  �D$ P�  �t$ ���L$Q����  �L$�:  _��^��� �ly�P�D$P�D$PQ�R$��� �����ly�P�D$P�D$PQ�R(��� �����ly�P�D$P�D$PQ�R ��� �����ly�P�D$P�D$PQ�R<��� �����ly�P�D$P�D$PQ�R,��� �����ly�P�D$P�D$PQ�R0��� �����ly�PDQ�R��ály�PDQ�R(��ály�PX�D$PQ�R8��� ����������ly�PX�D$PQ�R(��� ����������ly�T$�HDj j R���Ð���������ly�T$�HD�D$Rj P���Ð������T$�ly�HDRj h'  ���Ð�������Vj ��h�  �   �D$��tjj h�  ����   ����u^��� �L$�r����D$ Ph�  �L$�/����L$$Qh�  �L$�\����ly�B@j �L$QV�Pd���L$�����   ^��� �ly�PHj Q�Rd��Ð��������������ly�PH�D$P�D$PQ���   ��� ��ly�PH�D$P�D$PQ���   ��� ��D$VWP������������t�L$QV������_��^� ������D$VW���L$PQ����������t�T$RV���g���_��^� �ly�PH�D$P�D$PQ��(  ��� ��ly�HH�T$�D$R�T$P�D$R�T$PR���  ��Ð�����ly�T$�HHj R���Ð����������Vh�  �����������u^ËD$�L$PQ���i�����u�ly�B@V�PH��3���^Ð���������������ly�H@V�t$�R�QH���    ^Ð��ly�PHQ��8  ��Ð�������������ly�PHQ��$  ��Ð�������������ly�PHQ��(  ��Ð�������������D$�ly� Ð����ly���   �� Q���   YÐ����������VW�L$������D$$���|$ t%�ly�Q4P�R����u6�L$�9���_3�^��Ëly�B0W�P����u�L$����_3�^��Ë�L$Q�L$,Q���R$�L$���0������t�ly�B0�L$QW���   ���L$�����_��^��Ð�SVW�|$��������=ckhc��   ��   =TCAbatB=$'  t(=MicM�:  j hIicM���F����WP���R_^[� �W���P_^�   [� j hdiem�������WP���R_^[� =INIbt=NIVb��   ����P_^[� �F��t_^�   [� ����F   �R_^[� ����P_^[� =ytsddtL=ndmct(=dmmc��   �Wj hidmc������P���S_^[� �Wj hidmc���l���P���S_^[� ����R _�F    ^3�[� =atnit$=cnysu"j hIicM���.����WP���R_^[� ��  _^3�[� ��V����"�ly�H0Vh�G��F���F    ��^Ð�����V���   �D$t	V��	  ����^� ��V��F����"t�ly�Q0P�R���F    ^Ð������V��F��u^� �ly�Q0�L$ j j j j j Q�L$$j QjP���   �ly�B0�L$D�T$@Q�L$@R�T$@Q�L$<R�Vj QR���   ��D^� ������A��uËly�Q0P�R��Ð�������A����Vu�t$P���  ��^��� �L$�Q�	�5ly�v0R�T$RQP�D$P���   �t$$��P���  �L$�C  ��^��� �����������Q��u3�� �D$�H� V�5ly�v0Q�L$QPR�V��^� ����������������D$3҅���P�D$j BR�T$j PR�   � ��������������V��htniv�L$������D$(Phulav�L$����hgnlfhtmrf�L$�����L$,Qhinim�L$�s����T$0Rhixam�L$�`����D$4Phpets�L$�M����L$8Qhsirt�L$�:����D$$�T$RP�L$Q���������-  �L$���  �L$������^��� �Q��u3�� �D$�H� V�5ly�v0Q�L$QPR�V8�L$3҃��ɋL$��^�� ���������������Q��u3�� �D$�H� V�5ly�v0Q�L$QPR�V8��^� ����������������lyV�t$�VW���H4R��D$�F    �~�H� �ly�R0Q�L$QVP�GP���   ��3Ʌ����F_^��� ���������D$��u��y� �ly�I�R0V�t$VP�D$PQ�RP��^� ���������������ly�P0�Aj j j j j j j j j P���   ��(Ð��������   Ð����������   � ��������� �������������V�������#�F   �F    ��^�V���   �D$t	V�  ����^� ���#�����������D$�T$Vj P�D$��L$QRPj j ���������t�F��t	�   ^� 3�^� ���D$�A����� �S�\$V�������=ckhc��   tq=cksatW=TCAb��   Wj hdiem����������SW���F   �P�؋F��t��t��u3Ƀ���Q���~���_^��[� �F��tH����R^[� �F��t5���e�����t*�F    ^�   [� =atnit�D$PS�������^[� ^3�[� ��3�� @#�H�H�HÐ�����������V���   �D$t	V�K  ����^� ��V��FW3�;��@#u�ly�V�H4R����~�~_^Ð���ly�P4�AP�R��Ð�������������ly�P4�AP�R��Ð�������������ly�P4�D$�IP�D$P�D$P�D$PQ�R��� ��������ly�P4�D$�IPQ�R$��� �������ly�P4�D$(P�D$(P�D$(P�D$(�IP�D$(P�D$(P�D$(P�D$(P�D$(P�D$(PQ�RX��,�( ���������V��h�  �����D$�L$�T$P�D$QRP���8���^� ����QSVW�|$���3��=���=INIb��   ��   =SACb{t1=$'  t=MicM�I  _^��[Y� �W���P _�   ^��[Y� ��D$P�L$Q�Ή\$�\$�R��t�ly�L$�B4�T$Q�NRQ�P��_�   ^��[Y� =ARDb��   USj���$���j j�ϋ�����j j�ϋ��
���j j�ωD$ ������P�D$PSU���R]_�   ^��[Y� ����R_�   ^��[Y� =NIVbYtB=NPIbt,=ISIbuP�>�������P������P���W_�   ^��[Y� �W���P_^[Y� ����R_�   ^��[Y� =cnyst	_^��[Y� ShIicM���K����WP���R_^[Y� ������������D$j0P�t  ��ËD$j$P�d  �������@Ð��������ly�H�!�������ly�HV�t$�R�Q���    ^Ð��ly�P�D$P�D$P�D$PQ�R ��� ���������������V�t$���t�ly�QP�R���    ^Ð�������������D$�L$%�   S�؊���W�|$������f���ʃ��_[ËD$��s�   �ly�Qj j P��H  ��Ð����������D$��s�   �ly�Q�L$Q�L$QP��H  ��Ð����D$��t�ly�QP�RYÐ��������j�   ����u��`���������������D$hpyPh� ��  ��Ð�������V�t$�> t%j���������t��T$R�L$�P���    ^Ð��������������Vj����������t�@��t�L$�T$QR����^� 3�^� Vj���f�������t�@��t�L$�T$Q�L$RQ����^� 3�^� �����������Vj$���&�������t�@$��t�L$�T$QR����^� 3�^� VjH�����������t#�@H��t�L$�T$Q�L$R�T$QR����^� 3�^� ������VjT����������t#�@T��t�L$�T$Q�L$R�T$QR����^� 3�^� ��������3ɉ�H�H�H��   �����������V����t	P�������F���    t	P��������F    �F    �F    ^Ð�D$htyPh_� �  ��Ð�������VjH�����������t�@H��t	�L$Q����^� �����������VjT����������t�@T��t����^Ð�Vh�   ����������t0���   ��t&�L$�T$Q�L$R�T$Q�L$R�T$QR����^� ���^� ������Q3���~V�1���   @u	�����t@��Ju�^Ð���������lyV��HV�Q`����^Ð����������lyV��HV�Q`�ly�L$�BVQ�Pp����^� �������lyV��HV�Q`�L$�ly�Bj j�QV�Pd����^� ���ly�PQ�RlYÐ��ly�P�D$PQ�Rp��� ����������ly�T$V��HVR�Qp����^� ���V�t$���t�ly�QP�R���    ^Ð�������������ly�PQ�R��ËD$�L$��VPQ�L$��������"   �t$P��������L$�=�����^��Ð������D$V��P����P���K   ��^� ������D$P�   ���@� ���������������ly�P�D$j PQ�R ��� ��������ly�P�D$P�D$PQ�R0��� �����ly�P�D$P�D$P�D$PQ�RT��� ����������������ly�T$�HR�Q0YÐ��������������ly�T$�H�D$RP�QD��Ð�������ly�H�T$�D$R�T$P�D$R�T$PRh�#  ���   ��ály�T$�HR�QYÐ��������������ly�H�ap������ly�H�at������ly�H�ax������ly�T$�HR�Q|YÐ��������������ly�T$�HR���   YÐ�����������ly�T$�HR���  YÐ�����������ly�T$�H�D$RP���  ��Ð����ly�T$�H�D$R�T$PR���   ��Ð���������������ly�T$�H�D$R�T$PR��   ��Ð���������������ly�T$�H�D$RP��,  ��Ð����ly�P���D$ P�D$P�D$PQ��D  �L$���#���Ð���     �@    Ë��L$�    �H� �����������������L$�    �H� ���������������T$V���    �F    �ly���   j RV�Q����^� ��ly���   Q�Yály���   Q�R8��Ð�������������ly���   Q�R<YÐ��������������j�)   ����t�@��t�L$�T$Q�L$RQ�Ѓ��3�Ð���D$h�yPhD �<  ��Ð�������Vj\�����������t�@\��tV�ЋD$��P���&   ��^� Vj`����������t�@`��tV�Ѓ�^�Vjd����������t�@d��t�L$QV�Ѓ�^� ����������   �����������3��xy�|y��yÐ��������������ly���   �D$P�D$P�D$P�R� �ly���   �D$P�D$P�D$P�R � ��V��L$�q����ly�H �T$RV�Q �t$$���D$P�������L$�������^��� ������������ly�P �D$PQ�R$��� ����������ly�H\�!�������ly�H\V�t$�R�Q���    ^Ð��ly�P\�D$PQ�R��� ����������ly�P\�D$P�D$P�D$PQ�R,��� ����������������ly�H$�a������ly�T$�H$R�QYÐ��������������lyV��H$V�QD����^Ð����������lyV��H$V�QD�L$�ly�B$QV�P����^� �������lyV��H$V�QD�ly�L$�B$VQ�PL����^� �������ly�P$Q�RHYÐ��ly�P$�D$P�D$P�D$PQ�R��� �����������������V��L$�����ly�H$V�Q�����D$t�T$R���~����D$P�������t$�L$Q��������L$�H�����^��� ����������������� V��L$������ly�H$V�Q �����D$t
P�L$�   �T$R�  �t$,���D$P��������L$�������^�� � ��� V��L$�a����ly�H$V�Q$�����D$t
P�L$��   �T$R�&  �t$,���D$P���s����L$������^�� � ���V�t$$V�D$P�����������L$�m�����^��� �����ly�P$�D$PQ�R,��� ����������ly�P$�D$PQ�R0��� ����������ly�P$�D$PQ�R8��� ����������ly�T$V��H$VR�QL����^� ����D$��VP�L$�����ly�D$,�Q$P�L$Q�R@�t$,���T$R���u����L$������^��Ð����V�t$���t�ly�Q$P�R���    ^Ð�������������ly�H(�!�������ly�H(V�t$�R�Q���    ^Ð��ly�P(�D$P�D$P�D$P�D$P�D$P�D$PQ�R��� �ly�P(Q�R��ály�P(�D$P�D$P�D$PQ�R��� ����������������ly�P(�D$P�D$PQ�R��� �����ly�P(�D$P�D$PQ�R��� �����ly�P(Q�R$��ály�P(Q�R(��Ã�,V�t$4Vh�y�L$�����P�L$�������������L$�/����L$������^��,Ð���������������ly�PT�D$P�D$PQ�R��� �����ly�HTj hG  ���Ð�����������ly�HL�a������ly�PLQ�R ��ály�PLQ�R$��ály�PL�D$P�D$P�D$PQ�R0��� ����������������ly�PL�D$P�D$P�D$P�D$PQ�R4��� �����������ly�PLQ�R<��ály�PL�D$P�D$P���   � �������V��L$������D$Ph�  �L$�>����ly�QL�D$Pj V�R���L$�.���^��� ���������V��L$�����D$Ph�  �L$������ly�QL�D$Pj V�R���L$�����^��� ��������ly�T$�HR���   YÐ�����������ly�H���   ����8SUVW���b�����3�;�u_^]3�[��8� �L$������L$LQ�D$h]  �L$�\$0�\$8�\$<�\$@�\$L�D$D   �\$H�l$,�D$4�����ly���   SSU���P����   ���������;���   �ly���   ���R(���D$$Ph�   �t$0����������   �L$D;�t}�ly���   S���   ;�tf�ly���   V���R<�ly���   �T$DR���   ��;�t�ly�H@V�QH��;����h����L$$������L$�_���_^��][��8� �ly�B@U�PH�ly���   �D$HP���   ���L$$�����L$����_^]3�[��8� ���������������   � ��������V�t$���������^� ����������������   U��$�   ��u��$�   �2���3�]�Ġ   �W3��p������D$��   SV��$�   P�L$(�����h=�L$�����P�L$D�����t$Wj��L$,Q�T$LR��$�   P������P��$�   Q�������P�T$lR�������P���!�����K��ۍL$\�������L$x������$�   �����L$@�����L$�h����L$$����^��[t0��$�   �L$��$�   UP��$�   Q��$�   RPQ�>   �����T$R��������$�   �D$    ������_]�Ġ   Ð���������������   V��$�   ��u
3�^���   �j �D$h�   P������$�   ��$�   ��$�   h�   �L$T�L$Q�T$\��$�   �D$��$�   RPj�t$D�D$( i�D$l�h�D$p�h�D$t�h�D$x�h�D$|�h������ ^���   Ð���`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�� h#Ð�������h#Ð����������t�j�Ð�����D$��u��y�L$P�D$PQ�������Ð����������������3ɉ�H�H�H��   �����������V��F��Wu:���t�ly�Q<P�R���    �~��t���[���W�������F    _^Ð���������V�D$P���������P���   �L$��������^��Ð��V��F��W�|$u*j j j�F�������t
W�������3����Fu_^� �F��t�3���_��^� �ly�H<W���3҅��_�F   ^��� ����������������u�ly�H�� �ly�J<�T$RP�Q��� ������   �   ��������y����������h�j�  YÐ�����y������������y�����������D$P��y�q����V���l#�F    �ly�H4���   �F��^Ð����������V���   �D$t	V��������^� ��V��V�l#�ly�H4R���   3����F�F^Ð��������ly�P4�AP���   YÐ������������L$��t(�T$ �R�T$ R�T$ R�T$ R�T$ R�T$R�T$R�PÐ���������������D$�@�ly�R4V�t$Qh�kVP�AP���   ��^� ��V��������V�t#�ly�H4R���   �ly�H4�����   �F��^Ð�������V���   �D$t	V���������^� ���t#�����������ly�P4�D$�IP�D$PQ���   ��� ���������������ly�P4�D$�IP�D$PQ���   ��� ���������������ly�P4�D$�IP�D$PQ���   ��� ���������������ly�P4�D$�IPQ���   ��� ���� ��������������ly�P4�D$�IPQ���   ��� ����ly�P4�D$�IP�D$PQ���   ��� ���������������   � ��������� �������������3�� �����������3�� ������������   � ���������   � ���������D$�L$�T$�H4�L$�P �T$��L$�@ i�@8�h�@<�h�@@�h�@D�h�@H�n�@L�h�@P�n�@h�n�@X�n�@\�n�@`�n�@d�n�@Tpn�P0�H(�@,    Ë�`����������̋�` ����������̋�`$����������̋�`(����������̋�`,����������̋�`0����������̋�`4����������̋�`�����������3�� �����������3�� �������������   W3��������D$��   ��$�   SVP�L$$�S���h=�L$�U���P�L$@�;����t$Wj��L$(Q�T$HR��$�   P������P��$�   Q������P�T$hR�~�����P��������K��ۍL$X���A����L$t�8�����$�   �,����L$<�#����L$������L$ ����^��[t@��$�   �L$��$�   WP��$�   Q��$�   R��$�   P��$�   QRP�    �� ���L$Q��������_�Ġ   Ð�����   V��$8  W�����������$,  tj VW��������u	_^��   �j �D$h   P�%�����$T  ��$L  ��$P  Q��$D  R��$L  PQR�D$(P�3   ��$T  h   �L$0QRWj
������8_^��   Ð�������������D$�L$�T$V�t$P�D$Q�L$RPQV�������ǆ�   �qǆ�   Pqǆ�   `qǆ�   pq^Ð����������������`<����������̋�`@����������̋�`D����������̋�`8�����������V�t$��t���u9�D$jP�E�������u^Ë��U�����u^Å�t��p�T$3�;���I#�^Ð������D$H����   �$��r�   á�}@����}uL�L$Q������=L  }�����ËD$��u�����ÊV3���t��y+Ј�HF@��u�Ɔ�y ^�   ËT$�D$RP�����������H��3�����}u
�f����A����   Ã��ÍI �qxr}r�q�r]r�������������   ��  ��}�n  ���øk|��>y��>��>{y��>�x��>cy��>�U��� �EV�E�E��E�E�B   P�E��u�E����P�
  ���M��x�E��  ��E�Pj �	  YY��^��U��� �E�E�I   P�E�E��B  �E�EP�E��uP�r  �������������̋L$W��tzVS�ًt$��   �|$u��uo�!�F�GIt%��t)��   u����uQ��t�F�G��t/Ku�D$[^_���   t�GI��   ��   u����ul�GKu�[^�D$_É��It�����~�Ѓ��3��� �tބ�t,��t��  � t��   �uƉ�����  �����   ��3҉��3�It
3����Iu���u��D$[^_�U��� SV�uW�  j�EY3��}�j�_���ʋ�#�����D�F��u�U��u�E�P�j����[#������L5���t��tB���ڊ��t����j#�X�����L5���uB���" B�E_^�P��+����#�[����U������}��f�E���f�E��m��}��m��E�U��������Q=   �L$r��   -   �=   s�+ȋą���@PËD$����   � j��}��%  ��Yt<��}3Ɋ�}%�   �-�}��}��}�����}�E  ��u	� &  3��r�  �����"  ��}��  �   ��  �  ��}�>3�;�u,9�}~���}9�}u�  �G  �0  �%  ���uQ�  YjX� U��S�]V�uW�}��u	�=�} �&��t��u"�����t	WVS�Ѕ�tWVS�������u3��NWVS�������Eu��u7WPS�������t��u&WVS������u!E�} t�����tWVS�ЉE�E_^[]� ��}��t��u�=�}u�v%  �t$�%  h�   �@>YY�V�k  �5���{0  ���Y�����+��;�s=R�]0  ��P�5���-  ����u3��,���+�������������D$�������   ��^��t$�y������Y��H�h�   ��0  ��Y���uj�"������Y�  ���������������̺P>�a2  �P>��1  �Ƀ=�}t����@  �����z����h   h   �C  YY�U�����#�]���#�]��E��u��M��m��]��E��p!���vjX��3���h�#� ��th�#P� ��tj �������V�t$�P��D  ��eYt,F�=@B~�jP�MD  YY���LB�A����uԊDB��F�����F��u�^ËD$�DB���t:�t�H@��u�@��t*���t��et��Et@���H�80t�8uH�@A�҈u�ËD$� �#���rjX�3��U��QQ�} �ut�E�P��H  �EYY�M���M��H�ÍEP��H  �EYY�M���U���(�E�VP�E�P�EQQ� �$�lI  �u�E�P�U�FP3��}�-��3Ʌ�����Q��H  �E�j P�uV�u�	   �E��0^��U��S3�8]V�uW�}t3�9]��P3��>-���P�v  YY�>-��u�-�G9]~�P�H����DB�3�8]h�#���MQ��I  9]YY��t�E�FA�80t<�^Ky���-A��d|��jd�^�� �Ù����A��
|��j
�^�� �Ù���� Y��_^[]�U���(�E�VP�E�P�EQQ� �$�IH  �u�E�P�E��P3��}�-��EP�G  �E�j PV�u�	   �E��,^��U��SV�u�]W�FH�} t;Eu3Ƀ>-���ˋ�� 0�` �>-��u�-�{�F��jW�?  Y�0YG���} ~DjW�'  �DBY��vGY��}+�} t�����9u|�u�uW��   �uj0W�I  ��_��^[]�U���(SV�E�WP�E�P�EQQ� �$�KG  �E�]�p�3��}�-��E���E�PSW�F  �E��H;������|&;�}"��t
�G��u� G��E�jPS�u���������E�jP�uS�u������_^[��U��}et2�}Et,�}fu�u�u�u�N�����]��u�u�u�u�4�����u�u�u�u������]�W�|$��tV�t$V��  @PV�V��H  ��^_�U��SV�u�F�^����   �@��   �t�f ���   �N$���F�F�f �e $�f��Fu"���Dt���DuS�N  ��YuV�dN  Yf�FWtg�F�>+��H��NI���N~WPS�KL  ���E�6���t�ˋ����������������>�@ tjj S�8K  ���F�M��j�E_WPS��K  ���E9}_t�N ��E%�   � �F���^[]�U���H  SVW�}3��G�ۉu�u�}��  �M�3���M��u�3�9U���  �� |��x�Ê��#���3�����#�����E���  �$���M���ỦU؉U��U�U��U��x  �Ã� t;��t-��tHHt���Y  �M��P  �M��G  �M��>  �M���5  �M��,  ��*u#�EP��  ��Y�E��  �M��؉E��  �E��ˍ��DA���U���  ��*u�EP�  ��Y�E���  �M����  ���ˍDAЉE��  ��It.��ht ��lt��w��  �M��  �M��  �M� �  �?6u�4uGG�M���}�l  �UЋLB�U����DA�t�E�P�u��P�  ���G�}�E�P�u��P�f  ���%  �Ã�g�  ��e��   ��X��   �x  ��C��   HHtpHHtl����  f�E�0u�M��u����u�����EP�  f�E�Y�ȉM���  ��u	��>�M��E�   ����N����  f�8 ��  @@���E�   �� �M�@������;ʉ}���   �E�   ��   f�E�0u�M�f�E��EPt;�0  P������P�L  ���E��}2�E�   �)��Zt2��	t�H��  �  ��  Y�������E�   �������E���  �EP�  ��Yt3�H��t,�E�t� ��M��E��E�   �  �e� �M�� �  ��>�E�P�   u��gu�E�   �E�ũ��E�u��H��M��@��E���P������P�E�P��>�u�����   t�}� u������P��>Y��gu��u������P��>Y������-u�M��������}�W��  Y��  ��i��   ����   H��   HtQ�������HH��   ����  �E�'   �<+����  ��u	��>�M�����N��t�8 t@��+��  �E�   �E�   �E���E�   t]�E��E�0Q�E�   �E��H�E���E�   t;�M��5�EP�  �E� Yt	f�M�f���M��E�   �#  �M�@�E�
   �E��t�EP��  Y�A�E� t!�E�@�EPt��  Y����%�  Y�����E�@�EPt�  Y���  Y3��E�@t��|��s�؃� ���ڀM���������E��u�� �}� }	�E�   ��e�����u�e� �E��E��E��M������t;�E��RPWV�E��U��K  �uċ؃�0�u�WV�J  ��9����~]ԋE��M��뵍E�+E��E��E��E�t�M��90u��u�M�@�M��0�E�}� ��   �]���@t&��t�E�-���t�E�+�	��t�E� �E�   �u�+u�+u���u�E�P�uVj �  ���E�P�E��u�u�P�2  ����t��u�E�P�uVj0��   ���}� tA�}� ~;�E�]��x�f�CP�E�PC��H  Y��Y~2�M�Q�uP�E�P��   ����O��u���E�P�u�u��u��   ���E�t�E�P�uVj �q   ���}�G�ۉ}�����E�_^[�Øn~�~�~I�U��M�Ix��E�����Q�u����YY����Eu��]�� ]�VW�|$��O��~!�t$V�t$�t$�������>�t��O���_^�S�\$��KVW��~&�|$�t$�WF�t$P�u������?�t��K���_^[ËD$� � �@�ËD$� ��A��Q�ËD$� � f�@��U����  �e� SV�u3�W��]����]���	  �}��}3ۃ=@B~��jP��6  YY��LB���A��;�t6�M�W�E�WP�%
  YYP�
  �FFP��I  ����t�FFP��I  Y��>%��  �e� �e� �e� �e� �e� �e� 3��e� �]�]��]��E��]��^F�=@B~��jP�N6  YY��LB�ÊA����t�E��E����DCЉE��e��N>t^��*t2��FtT��It
��Lu7�E��E�~6u,�~4�Fu#�EЃe� �e� ���'�E��"��ht��lt
��wt�E���E��E���M��M��}� �O����}� �uu�E�E����E�@��EԀe� �}� u�<St
<Ct�M����E��]�3�� ��n�u�t(��ct��{t�u�E�P�  Y��u�E��v  Y�E�3�9E�t	9E���  ��o�^  �
  ��c�,  ��d��  �j  ��g~8��it��n�W  �}� �}��   �!  jd^�]��-�~  �E��z  �]썵<�����-u��<�����=������+u�}�M��E�W��  ��Y�]���}�}� t	�}�]  ~�E�]  �=@B~jS�n4  YY��LB�X����t!�E��M��t�E�F�E�W�p  ��Y�]��8DBuf�E��M��t\�E�W�M  �ؠDB�Y�]�F�=@B~jS� 4  YY��LB�X����t!�E��M��t�E�F�E�W�  ��Y�]�뻃}� ��   ��et	��E��   �E��M��tv�eF�E�W��  ��Y��-�]�u�F���+u�E��M��u!E���E�W�  ��Y�]�=@B~jS�Y3  YY��LB�X����t�E��M��t�E�F��M�WS�r  �}� YY��  �}� �M  �È& ��<���P�E��u�HP��>���)  9E�u
�E��E�   �}� ~�E���>�  �ƃ�p��  ����   HH��  ���������t$�;E��?  �M�}� ��  �E��E�  �}� ~�E��}G�}�?^��   �Ǎx�   ��+u"�M�u�}� t�E���u�E��h  ��Y�]��0�E  �u�E��N  ��Y��x�]�t/��Xt*��x�E�   tjo^�  �u�M�S�8  YYj0[��  �u�E��	  Y�؉]�jx�π}� ~�E���>�M��j �E�j P��9  ���}�{u�?]u	�]G�E� ��Uˊ<]t_G<-uA��t=���]t6G:�s�����:�w!����+�F�ʋ������D�BNu�2���ȊЋ��������D�뛀? �  �}�{u�}�}�u��M�W�u�u��S  YY�}� t�E��M����   �E�W�  ���Y�E�t~��j��Z�]�������L�3˅�t`�}� uR�}� tA�LB�E����DA�t�E�W��  Y�E��5@B�E�P�E�P�B  f�E�f�FF��F�u��d����E��\����M�WP�  YY9u��(  �}� �  �Ẽ}�c�r  �}� �E�t	f�  �`  �  �X  �E��]��-u�E����+u"�M�u�}� t�E���u�E��  Y�؉]�}� �  �}� ��   ��xuO�=@B~h�   S�/  YY��LB�X%�   ����   �E؋U�jY�1C  S�E؉U��}  ��Y�]��S�=@B~jS�m/  YY��LB�X����t]��ou��8}S�E؋U�jY��B  �j j
�u��u��B  �E؉U��E�CЙE�U܃}� t�M�t$�u�E��6  ��Y�]��+����u�M�S�9  YY�}� ��   �E؋M��؃� �E��ىM���   �}� ��   ��xt?��pt:�=@B~jS�.  YY��LB�X����tv��ou
��8}l���?�<����8�=@B~h�   S�k.  YY��LB�X%�   ��t7S���D  ��Y�]��E�}� �|�t�M�t$�u�E��X  ��Y�]��\����u�M�S�[  YY�}� t�߃�Fu�e� �}� ��   �}� u)�Ẽ}� t�EԋM؉�M܉H��}� �E�t�8�f�8�E��E�u�B�E�W��   ��Y�F;É]�uuU�LB���DA�t�E�W�   Y�F;ȉuu>�M��}��u�>%uM�E�xnuD������V����0�u�M��u���M�WS�   YY��M�WP�}   �M�WS�s   ���}��u�E̅�u8E�u�����E�_^[�Ã=@BV~�t$jV��,  YY��t$�LB�p����u��߃���^ËT$�Jx	�
�A�
�R�x@  YÃ|$�t�t$�t$�>A  YY�V�t$W�t$�������W�?  Y��Yu��_^������������̋L$��   t�A��t@��   u�    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��V�5B  � �����>t:jtj��@  ��Y��Yt)V�5�>� ��tV�4   Y� �N�j�X^�3�^��B  ��>���tP� ��>�ËD$�@P�G�@   �VW�( �5�>���$ ����u?jtj�T@  ��Y��Yt&V�5�>� ��tV����Y� �N���j�����YW�  ��_^á�>�����   V�t$��uP�$ ����tl�F$��tP�)B  Y�F(��tP�B  Y�F0��tP�B  Y�F8��tP��A  Y�F@��tP��A  Y�FD��tP��A  Y�FP=�GtP��A  YV��A  Yj �5�>� ^á0>��t��h 0h0��   h0h 0��   ���j j�t$�   ���jj j �   ���W�   j_9= ~u�t$�4 P�0 �|$ S�\$�=�}��}u<�����t"���V�q�;�r���t�Ѓ�;5��s�^h,0h$0�C   YYh40h00�2   YY��[t�   _��t$�= ~�, _�j�K@  Y�j�@  Y�V�t$;t$s���t�Ѓ���^�U���HSVWh�  ��  ��Y��uj����Y�5�����    ���  ;�s�f ���f �F
�����$�  �ލE�P�D f�}� ��   �E����   �8�X�;�E��   ;�|��9=��}V���h�  �6  ��Yt<��� ����  ;�s�` ���` �@
���$���  ����9=��|���=��3���~L�E�����t8��t2�uQ�@ ��t#�΋��������������M��	���H�E�FC;�|�3ۋ���ۃ<���4�uM���F�uj�X�
��H������P�< �����tW�@ ��t%�   �>��u�N@���u
�N��N�C��|��5���8 _^[��SVW������t7���  ;�s!�_�{� tS�H ���$�  ��$;�r��6�>  �& Y������|�_^[�S3�9��VWu�;C  �5�}3��:�t<=tGV����Y�t���   P�  ��Y;�5�}uj	�����Y�=�}8t9UW�f�����YE�?=t"U�Y  ;�Y�uj	����YW�6��-  Y��Y�8u�]�5�}��=  Y��}�_^���   [�U��QQS3�9��VWu�}B  �~h  VS�L ����5�}��8t���E�P�E�PSSW�M   �E��M���P�  ����;�uj�����Y�E�P�E�P�E���PVW�   �E���H�5�}_^��}[��U��M�ESV�! �uW�}�    �E��t�7���}�8"uD�P@��"t)��t%����a�t���t��F@���tՊ�F�����t�& F�8"uF@�C���t��F�@����a�t���t��F@�� t	��t	��	ū�uH���t�f� �e �8 ��   ��� t��	u@��8 ��   ��t�7���}�U��E   3ۀ8\u@C���8"u,��u%3�9}t�x"�Pu����}�}3�9U�U���K��tC��t�\F�Ku���tJ�} u
�� t?��	t:�} t.��t����a�t�F@���F�����a�t@��@�X�����t�& F�������t�' �E_^[� ]�QQ�SU�-` VW3�3�3�;�u3�Ջ�;�t�   �(�\ ��;���   �   �   ����   ;�u�Ջ�;���   f9��t@@f9u�@@f9u�+Ƌ=X ��SS@SSPVSS�D$4�׋�;�t2U�&  ;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$��:  Y�\$�\$V�T ���S��uL;�u�\ ��;�t<8��t
@8u�@8u�+�@��U�  ��Y;�u3��UWV�J?  ��W�P ���3�_^][YY�V�t$j �& � f�8MZu�H<��t��H��@�F^�U��,  �	�����h���SPǅh����   �h ��t��x���u��l���rjX�  ������h�  PhL$�d ����   3ۍ�����8�����t�<a|<z, �A8u퍅����jPh4$�E  ����u�������I��d���h  PS�L 8�d�����d���t�<a|<z, �A8u퍅d���P������P�HD  YY;�t>j,P�zC  Y;�Yt0@��8t�9;u��A8u�j
SP�A  ����t��t��t�E�P�����}�Y���[��3�j 9D$h   ��P�p �����t6���������uh�  �mD  Y�
��u�O  ��u�5���l 3��jXá��V��WufS3�90�U�-x ~@�4��=t �ph @  h   �6��h �  j �6���vj �5���Ճ�C;0�|��54�j �5����][�'��u"�PI���F��th �  j P�t �6;�u��5���l _^á�}��t��u*�=�}u!h�   �   �Y��t��h�   �   Y�U���  �U3ɸ ?;t��A=�?r�V����;� ?�  ��}����   ��u�=�}��   ���   ��   ��\���h  Pj �L ��u��\���h<'P��&  YY��\���WP��\����C���@Y��<v)��\���P�0�������\�����;j�h8'W���������`���h'P�&  ��`���WP�&  ��`���h'P�&  ��?��`���P�&  h  ��`���h�&P�XT  ��,_�&�E��?j P�6����YP�6j��< P�| ^��U��M3�SV�A�MWj�A�M[�A�M��t�E�E�  �	X��t�E�E�  ��H��t�E�E�  ��H��t�E�E�  ��H��t�E�E�  ��H�u�Ej��P��#˃�����_�H��E�ыP������ʉH��E�ыP������ʉH��E�ыP��#σ��ʉH��E�ыP��#˃��ʉH��  ��t�M�I�t�M�I�t�M�I�t�M	y� t�E	X��   #�t4=   t=   t;�u(�E�� �E������
�E����ˉ��E� ���   #�t =   t;�u"�E� ���E�������E�������E�M���  ����� ��ʉ�E	X �E�H ���ωH �E� �E�X�E	XP�E�HP���ϋ}�HP�E��X@��  �EPSj �u�� �E�@t�&��@t�&��@t�&��@t�&�Xt�&ߋ��������� t%ItIt	Iu�N����������������!������� tItIu!��#ʀ���#ʀ���@@�_^[]�U����ESW����j�[t�]tS�G  Y�����  �t�Etj�-  Y����  ����   �E��   j�  Y�   �M#���   ��   tX��   t(;���   �M��#�x@���w���]��E��n�M��#���v�h@��x@���]��E��F�M��#���v�x@��h@���]��E���M��#�h@���w���]��E�������   ���   �E��   V3��t��E� �]��E��#�����   �E�E�PQQ�$�  �E����]� ���������}	����]��T�E��#���s���3ҊE���f�E�����;�}+��]�t��u���m�]�t�M���m�Hu��t�E����]��E�E�����^tj�x  Y����Et�E tj �a  Y���3���_[���ËD$��t~���FP  � "   ��:P  � !   �U��QQ�E�M�E�  f����]����f�E��E���U��QQ�E�#V���u��3��]��   3�f�E�ue�E�� u9MtW�E�#�������sjX�3��Eu�e�E�t�M�eN��f�e��;�t�M��EQQQ�$�P����]����'�EQQQ�$�:����E���]���f%������  �E�E��0^��U��Q��}��E���U��Q�}����E���U��Q��}��E��#E��#M�ȉM�m�E���U��QQ�M��t
�-�@�]���t����-�@�]�������t
�-�@�]����t	�������؛�� t���]����U��j�h(h��d�    Pd�%    ��(SVW�]3�;�u�u��  Y��  �u;�uS�/  Y��  ������9  �}܃����   j	��.  Y�}�S�s;  Y�E�;���   ;58�wLVSP�`C  ����t�]��8V�>  Y�E�;�t*�C�H�E�;�r��PS�u���3  S� ;  �E�SP�A;  ��9}�uK;�uj^�u������uVW�5���� �E�;�t#�C�H�E�;�r��PS�u��3  S�u���:  ���M���Z   9}�u";�uj^������uVSW�5���� �E܋E�;���  9=���  V�SM  Y��������  �u�]3�j	�5.  YÃ��G  ���w;�v������j^�u�}܃����   j	�-  Y�E�   �E�P�E�PS�iG  �����}Ѕ���   ;5tis\����SW�u��u��K  ����t�E�E��8S��G  Y�E܅�t*����E�;�r��P�u�u��|2  W�u��u��RG  ���]�}� uSVj �5���� �E܅�t=����E�;�r��PS�u��52  W�u��u��G  ���VSj �5���� �E܃M���&   �E�;�uf9=�t^V� L  Y��������K�u�]j	��,  Y3��3����w;�uj^�����VSW�5���� ;�u9=�tV�K  Y��u�3��M�d�    _^[��U��j�h (h��d�    Pd�%    ��SVW�����uFj	�,  Y�e� �uV�z8  Y�E��t�v���	�u���u��M���	   �}� �U�u�j	�',  YÃ�uFj	�+  Y�E�   �E�P�E�P�u�E  ���E؅�t�0���u���u��M���-   �}� u�uj �5���� ���ƋM�d�    _^[�Ëu�j	�+  Y��5��t$�   YYÃ|$�w"�t$�   ��Yu9D$t�t$�uJ  ��Yu�3��U��j�h8(h��d�    Pd�%    ��SVW�����uC�u;58���   j	��*  Y�e� V�:  Y�E�M���   �E��tm�   j	��*  YÃ�uZ�E��t�p����j^�u;5tiw.j	�r*  Y�E�   ����P��D  Y�E�M���   �E��u-V��uj	�*  YËE��ujX��$�Pj �5���� �M�d�    _^[������U���0���S�ٽ\�����=�j t�  ��8����   [����ݕz������U���U���0���S�ٽ\����=�j t�  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����  �   [�À�8�����=�} uLݕ0�����p���
�t<�t@<�t<
�t0����r����   f��\���f�� u���f�� tǅr���   �z٭\�����f��6���f%�f�tf=�t0�ǅr���   �h(�����������X(����s4�x(�,ǅr���   �`(�����������P(����v�p(VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�jI  ��_^�E��$���U���0���S�u�u�   ���ٽ\�����8�����J   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�������̀zuf��\���������?�f�?f��^���٭^�����@�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����@�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����@���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�@��p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t��������@ u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t��@����@���l$�����@����@���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ��������@�|$�l$�ɛ�l$������l$��Ã�,��?�$�>A����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������@ �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����,A�Ƀ�u�\$0�|$(���l$�-4A�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�A�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���A�|$�A�<$� �|$$�D$$   �D$(�l$(���A�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������@ �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����,A�Ƀ�u�\$0�|$(���l$�-4A�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�A�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���A�|$�A�<$� �|$$�D$$   �D$(�l$(���A�<$�l$$�Q�����0Z�����0Z�������@����������U��QV��}��u��:   ���E��#��E#E�V�   Y�EY�m��^�ËD$%����P�t$����YY�S�\$3�U��WtjX��t��t��t�� t��t   ��V�Ѿ   �   #ֽ   t��   t��   t;�u������#�^t;�u   �   _]��[t   �S�\$3�V��tjX��t��t��t��t ��   t�˺   #ʾ   t��   t;�t	;�u���������ˁ�   t��   u���^��   [t���U��Q�E�H��   w�LB�A�R��V�5LB�����DV�^t�e� �M��E�j�	�e� �E�jX�M
jj j QP�E�Pj�8  ����u���E
#E��S3�9�u�D$��A|Y��ZT�� [�V��WV�� 9��=� tV��j�!  Yj[�t$�   ��Y�D$t
j�e  Y�V�׋D$_^[�U��Q�=� SVWu�E��A��   ��Z��   �� �   �]�   j;�^}%95@B~VS�����YY�
�LB�X#ƅ�u���e�LB�������DJ�t�e
 j�E�]	X�	�e	 �]��Vj �M�jQP�EPW�5��8  �� ��t�;�u�E���E��M����_^[�ËD$Vj �Y��j���D$���Y�D$+ʃ�����҅�uF��}���8 uF����|�jX^�3�^ËD$SVWj �\$�Y�����D$����<�WjYjX+���P�7�g:  ��Nx�<���tWj�7�P:  ��N����}�_^[�U��QQ�ESVW�x�j Y�e� �_j ��^���j�ȋÙ���E^j�M����E+�Z����t!CS�u����Y��YuW�u�N���Y�E�Y�E�������jY!�E�@;�}�U+ȍ<�3��E�_^[�ËD$�L$Vj+�Z�0�4��Ju�^�W�|$3����_ËD$3Ƀ8 uA����|�jX�3��U����ESVWj �}[�������E�   ���E�E����e ����+��֋��#ΉM�����E��E��˃����M��Eu܋}�j[��jY��;�|�U��+Ƌ���E�$ K��y�_^[��U����ESVW�H
�ف� �  �M�H�M�H� �}���  ���?  �M���������E�u&�E�3�P������Y��   �E�P�����YjX��   �E�P�E�P�����w�E�P��������tC�G��+O;�}�E�P����Y�<;�?+Ë��E�P�E�P�v����E�VP�����w�E�P������G@P�E�P������ 3��|���;|(�E�P�V����w�M���E�P�m����w��7j�R����w�w�e��E�P��I���YY3�jY+O���M��Ɂ�   ��u��@u�M�U��q��
�� u�M�1_^[��hXD�t$�t$�������hpD�t$�t$�l������U���3�PPPP�u�EP�E�P��8  �u�E�P������$��U���3�PPPP�u�EP�E�P�8  �u�E�P������$��U��US�]V�u�JW�~�0�ۋ�~�]3ۊ��t��A�j0Z�@�Mu�U�  ��|�95|H�89u� 0��� �>1u�B�W����@PWV�u  ��_^[]�U���(V�EWP�E�P�G   Y�E�Y�u�Pj j������f��<  �u�}�F�Eډ�E؉F�E�PW��   �� �~��_^��U��Q�USVWf�B��  ��% �  ��#ωE�B��پ   �%�� �ۉu�t;�t�� <  �(��  �!3�;�u;�u�E�X�f�X�K��<  �]�������ȋEM����H���u�ɋ���ٍ��X����  ���ߋM�f�H_^[�������������W�|$�j��$    ���L$W��   t�A��t;��   u�����~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�A��td�G��   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_ËT$�L$��tG3��D$W����r-�ك�t+шGIu������������ʃ���t��t�GJu��D$_ËD$���������U��WV�u�M�}�����;�v;��x  ��   u������r)��$����Ǻ   ��r����$���$����$���� �L�p�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ�F��G��r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������0��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�@��I �Ǻ   ��r��+��$����$�����������F#шGN��O��r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������Z�������$����I D�L�T�\�d�l�t����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��j�)���Y�V�t$;5��s@�΋������������D�t%WV�i:  �t$�t$V�(   V���:  ����_^��*  � 	   �*  �  ���^�V�t$WV��9  ���Yu��)  � 	   �-�t$j �t$P�� �����u�( �3���tP�G)  Y�����΃����Ƌ������d���D���_^�V�t$;5��s@�΋������������D�t%WV�9  �t$�t$V�(   V����9  ����_^��@)  � 	   �>)  �  ���^�U���  SVW3�9}�}��}�u3��f  �E�������E���4�����D0 tjW�u����������@���   �E9}�E��}��   �������M�+M;Ms)�M��E��	��
u�E�� @�@�ȍ�����+ʁ�   |̋�������+��E�j P������WP��40�| ��tC�E�E�;�|�E�+E;Er�3��E�;���   9}tbj^9uuL�((  � 	   �&(  �0�A�( �E�ǍM�WQ�u�u�0�| ��t�E�}�E���( �E��u�f'  Y����,��D0@t�E�8������'  �    �'  �8��+E�_^[���h   �����Y�L$���At�I�A   ��I�A�A�A   �A�a �ËD$;��r3�Ëȃ����������D���@á��Vj��^u�   �;�}�ƣ��jP��  Y�h���Yu!jV�5����  Y�h���Yuj蠪��Y3ɸ�D�h���� ��=G|�3ɺ�D��������4����������t��u�
��� A�� E|�^��B8  �=�} t�)7  ËD$��D;�r=�Fw+�����P�
  YÃ� P�� ËD$��}��P��  YËD$�� P�� ËD$��D;�r=�Fw+�����P�  YÃ� P�� ËD$��}��P��  YËD$�� P�� �U��SV��WV�� �=� 3�9�tV��j�\  Yj[�u�u�   Y�E��Yt
j�  Y�V�׋E_^[]�U��E��u]Ã=� uf�Mf��� w9j�X]ÍM�e Qj �5@BP�EjPh   �5��X ��t�} t�%  � *   ���]������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� U��SV��WV�� �=� 3�9�tV��j�  Yj[�u�u�u�   ���E��t
j��  Y�V�׋E_^[]�U��SV�u3�;�t9]t�:�u�E;�tf�3�^[]�9�u�M;�tf��f�jX��LB���DA�tN�@B��~*9E|/3�9]��Q�uPVj	�5��� ���@Bu�9Er8^u��/#  � *   ����3�9]��P�ujVj	�5��� ���x����Ƀ=@B~j�t$�����YYËD$�LB�A���������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̀�@s�� s����Ë�3������3�3��V�t$�F����   �@��   �t
 �F�   f��Fu	V����Y��F��v�v�v�4  ���F��to���tj�V�u7�NW���t�������<����ɍ<����>�O_�ႀ��u�� �V�~   u�N��t��u�F   �H�F�A�^��������	F�f ���^�S�\$���VtA�t$�F�u��t2�u.�~ uV�����Y�;Fu	�~ u@��F@t��8t@����^[�����F�F$��F��%�   ��U��j�h�(h��d�    Pd�%    ��SVW�u�u�u�u���w3�;�uj^������u�3ۉ]������   �����uA�}�;=8�w|j	�_  Y�]�W�.  Y�E��M���   9]�t^�u��H3ۋuj	�  YÃ�uA;5tiw9j	�  Y�E�   ����P�  Y�E��M���L   9]�tVS�u��2�����9]�u>Vj�5���� �E�9]�u'9�tV�"   Y���0����3ۋuj	�
  YËE��M�d�    _^[��V�5� �5TG���5DG���54G���5G��^�VW�=H �G���t+��TGt#��DGt��4Gt��GtP���6�   Y�����G|��54G���5DG���5TG���5G��_^�U��EV�<�G �4�Gu>Wj������Y��uj�ܢ��Yj������> YWu
�� �>��*   Yj�   Y_�6�� ^]�U��E�4�G�� ]�U��j�h�(h��d�    Pd�%    ��SVW�u����   �����u;j	�K���Y�e� V��  Y�E��t	VP��  YY�M���   �}� �Qj	�z���YÃ�uSj	����Y�E�   �E�P�E�PV��  ���E܅�tP�u��u��  ���M���   �}� u�u�
j	�"���Y�Vj �5���x �M�d�    _^[��U���SVWj�����u�  ��Y;<�Y�]u3��p  ���V  3Ҹ`H9tt��0B=PIr�E�PS�� j^;��!  j@�%d� Y3��`�9u�󫪉<���   �}� ��   �M�����   �A���;���   ��a�@��e� j@Y3��`��4R������pH�; ��t,�Q��t%���;�w�U���XH�a�@;�v�AA�9 u��E����}�r��E�L�   P�<���   ��dH�@���Y�d���RAA�y� �G����ƀ�a�@=�   r�S�   Y�d��5L���%L� 3��@������=x t�   �   �������j�]���Y��_^[�ËD$�%x ���u�x   �%� ���u�x   �%� ���u���x   ËD$-�  t"��t��tHt3�ø  ø  ø  ø  �Wj@Y3��`��3��@��<��L��d����_�U���  �E�VP�5<��� ���  3��   ������@;�r�E�ƅ���� ��t7SW�U��
��;�w+ȍ�����A�    �����˃��BB�B���u�_[j �������5d��5<�P������VPj��  j �������5<�VP������VPV�5d���  j �������5<�VP������VPh   �5d���  ��\3�������f���t��a���������`����t��a� �������〠`� @AA;�r��I3��   ��Ar��Zw��a��Ȁ� ��`����ar��zw��a� �Ȁ� ����`� @;�r�^�Ã=�� uj�����Y���   ���U��WV�u�M�}�����;�v;��x  ��   u������r)��$����Ǻ   ��r����$����$�����$�<������ �#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ�F��G��r���$����I ������|�t�l�d�\��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�@������$����I �Ǻ   ��r��+��$�H��$�@��X�x����F#шGN��O��r�����$�@��I �F#шG�F���G������r�����$�@���F#шG�F�G�F���G�������Z�������$�@��I ��������$�7��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�@���P�X�h�|��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��j �t$�t$�t$�   ���U���S�e� VW�}��w�u��=@B~��jP�Y���YY��LB�ÊA����t�F�Ѐ�-�u�u�M���+u�F�u��E����  ����  ��$�w  j��Yu$��0t	�E
   �2�<xt<Xt	�E   ��M9Mu��0u�<xt<Xu�^FF�u����3��u�  �E�=@B��~jV����YY��LB�p����t�˃�0�2�=@B~WV�q���YY��LBf�p#ǅ�tJ��P�!*  Y�ȃ�7;Ms6�u��M;u�ru���3��u;�v�M�	�u�u��E��E���d����E�M��]�u��t�E�E��e� �K�����u�u>��t	�}�   �w	��u,9u�v'��  �E� "   t�M����E$�����ƉE���t�E���Et�E��؉E��E���E��t�83�_^[����������������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
B8�tф�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[����̋L$WSV��|$��ti�q��tO���L$�F8�t��t�F8�t
��u�^[_3�ÊF8�u�~��a��t(���8�uĊA��t�f���8�t��3�^[_��������G�^[_Ë�^[_�U��WVS�M�&�ً}��3����ˋ��u�F�3�:G�wtII�ы�[^_��h@  j �5���� ���4�uËL$�%,� �%0� j�(��8�� �   Xá0����4���;�s�T$+P��   r����3��U����MSV�u�AW�����+y����i�  ��D  �M��I���M���  �1�1�U�V��U��U����]u~��J��?vj?Z�K;KuL�� s�   �����L��!\�D�	u(�M!�!�J�   ���L��!���   �	u�M!Y�M��]��M��S�[M�Z�U�M��Z�R�S����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M��щM���J;�v��;�tc�M�q;qu@�� s�   �������!t�D�Lu&�M!1��K�   �����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��\��щ^�N�q�N�q�N;Nu`�L�� �M���Ls%�} u�   �����M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �,�����   �$��5t ��H� �  h @  SQ�֋$��,��   ���	P�,��$��@����    �,��@�HC�,��H�yC u	�`��,��x�uiSj �p�֡,��pj �5���x �0��4������ȡ,�+ȍL�Q�HQP�����E���0�;,�v�m�4��(��E�=$��,�_^[��U����0��4�SV��W�<��E�}��H����M���I�� }�����M���u��������3���u�E��(���;߉]s�K�;#M�#��u��;]��]r�;]�uy��;؉]s�K�;#M�#��u����;�uY;]�s�{ u���]��;]�u&��;؉]s�{ u����;�u�8  �؅ۉ]tS��  Y�K��C�8�u3��  �(��C�����U�t����   �|�D#M�#��u7���   �pD#U�#u�e� �HD֋u�u���   �E�#U�����#9�t�U���3�i�  ��D  �M�L�D#�u����   j #M�_��|��G���M�T��
+M���M���N��?~j?^;��  �J;Jua�� }+�   �����M��|8�Ӊ]�#\�D�\�D�u8�]�M�!�1�O�   ���M��|8����   ��!��]�u�]�M�!K��]�J�z�}� �y�J�z�y��   �M�|���z�J�Q�J�Q�J;Jud�L�� �M})���} �Lu�   �����	;�   �����M�	|�D�/���} �Lu�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;,�u�M�;$�u�%,� �M���B_^[�á0�� �VW3�;�u0�D�P��P�54�W�5���� ;�ta� ��4��0��4�h�A  j���5���4��� ;ǉFt*jh    h   W�� ;ǉFu�vW�5���x 3���N��>�~�0��F����_^�U��Q�MSVW�q�A3ۅ�|��C����j?i�  Z��0D  �E��@�@��Ju��j��yh   h �  W�� ��u����   �� p  ;�w<�G�H�����  ����  �@��  ��������Hǀ�  �     �H�;�vǋE��O�  j_�H�A�J�H�A�d�D ����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ESVW�}�׍p+Q�A�������i�  ��D  �M�O�I;�M�\9��|9��]��_  ���O  �;��E  �M���I��?�M�vj?Y�M��_;_uH�� s�   ���M��L��!\�D�	u+�M!�$���   ���M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;Yu\�L�� �M���Ls!�} u�   �����M	�D�D�   ����%�} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��G  3��C  �:  �])u�N�K��\3��u�]��N�K���?vj?^�E���   �u���N��?vj?^�O;OuG�� s�   �����t��!\�D�u(�M!�!�N�   ���L��!���   �	u�M!Y�]�O�w�q�O�w�q�uu��u��N��?vj?^�M�|���{�K�Y�K�Y�K;Ku\�L�� �M���Ls!�} u�   �����M	9�D�D�   ����%�} u�N�   ���M	y����   �N�   ���	�E��D�jX_^[�Ã=`I�SUVWu�PI�h    j �5���� �����  �-� jh    h  @ j �Ջ�����   j�   h   SW�Յ���   �PI;�u�=PI u�PI�=TI u�TI���TI�F�5TI�F�0��  @ ���   �F�F�N�~�F3��   3҃���J#�JE��H����   |�Sj W��������F�;�s���   ��G��G�   ��   �܋��'h �  j W�t ��PItVj �5���x 3�_^][�V�t$h �  j �v�t 95piu�F�pi��PIt �F�Vj ���N�H�5���x ^Ã`I�^�U��QSV�5TIW�~���   �e� ��   � �? �?�   u9��h @  Fh   P�t ��t���|�F��t;�v�~�E��Mt��   ����}��}� �΋vt,�y�u&j�A Z�8�uB����   |��   uQ� ���Y;5TIt
�} �P���_^[�ËD$�PIV��;Av;Ar�	;�t7��u1��   ���  ;�r �t$��t$��f�� �+��+�^���D�3�^ËD$�L$+H���D��L$��! �8�   �@�   u�|�=| uj����Y�U��QQSV�5piW�V�����   �~��   ��+ƃ������;��E�s:��];�|9_vSQP�  ����uu�E��_����      ;��E�r���]�F�N�~�E�;��M�s3�;�|9_vSP�u��j  ����u&�_�E�   ��;}�r���]�6;5pit�C����5pi)�~�(  �PI����t� u�?;���   ��_�e� ���+�������w�;�u�}�}���E��8�t�E�j��h   PV�E��� ;���   j �u�V�u����U����ҋ�~0�F�U����   ��P�P���   ���A�      ���M�u։=pi��   ;�s�9�t����;��#��G�E�F�_))F�L��   ��4�4�����t)�H�Y�T�pi���   +ӉQ��)P��   �3�_^[��U��Q�M�USV�qW�9���   ;�}��ǉ]r!��;�s)Q�	�a �A��G��   ��> t�ƍ4;�sC���u0j�X^�; uCF��;�sN;E�u�q�)u9U��   �}������ƍ4;ur��q;�s~�;Esv���u@j�^X�; u%C@���;]s	+��q�	�a �q�1����6;�s)E9Ur4������맍;]s	+�A�	�a �A���Fk���+��3�_^[��U��Q�US�]V�
W�}�e� ��+G��;M�|�v�E+Ȉ�G�   �`se�E�4���   ;�wU�;�s
�8 u@��;�uB�E��;�w+;�v'���   ;�s3��38u@�< t��C�	�c �C�+M�E�   �E�_^[��S3�9�VWuBh�(�� ��;�tg�5 h�(W�օ���tPh�(W��h�(W���֣�����t�Ћ؅�t����tS�Ћ��t$�t$�t$S��_^[�3���V�v   �L$3���xi;t"��F=�jr��r"��$w�B   �    ^��5   ��|i^�Á��   r���   w�   �    ^��   �    ^��c�������Z������3�á���t�t$�Ѕ�YtjX�3��U��SVWUj j h���u�<  ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�h��d�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ��j�
SQ��j�M�K�C�kY[� ��VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{���ta�v�|� tEVU�k�T�]^�]�t3x<�{S�������kVS��������vj�D��a������C�T��{�v�4�롸    ��   �U�kj�S������]�   ]_^[��]�U�L$�)�AP�AP�y�����]� U���X�ESV�u��WH�Mt+Ht$HtHtHtHHtHunj��   �bj�
j�j�j[�~QWS�;�������uA�E��t��t��t�e����M��F����]Ѓ��M��NWQP�ESP�E�P�C�����h��  �u�,����>YYt�=�j uV�T�����Yu�6�۬��Y_^[��U��j�h�(h��d�    Pd�%    ��SVW�e表3�;�u>�E�Pj^Vh�(V�� ��t����E�PVh�(VS�� ����   jX����u$�E;�u���u�u�u�uP�� �   ����   9]u���ESS�u�u�E �����@P�u�� �E�;�tc�]��< �ǃ�$��d~���e��u�WSV�4������jXËe�3�3��M��;�t)�u�V�u�uj�u�� ;�t�uPV�u�� �3��e̋M�d�    _^[��U��j�h)h��d�    Pd�%    ��SVW�e�3�9=�uFWWj[Sh�(�   VW�� ��t���"WWSh�(VW�� ���"  ��   9}~�u�u�  YY�E����u�u�u�u�u�u�u�� ��   ����   9} u���E WW�u�u�E$�����@P�u �� �؉]�;���   �}����$���|���e�ĉE܃M���jXËe�3��}܃M���]�9}�tfS�u��u�uj�u �� ��tMWWS�u��u�u�� ���u�;�t2�Et@9}��   ;u�u�uS�u��u�u�� ����   3��eȋM�d�    _^[���E�   �6��$��I|���e�܉]��M���jXËe�3�3ۃM���u�;�t�VS�u��u��u�u�� ��t�9}WWuWW��u�uVSh   �u �X ��;��q������l����T$�D$��V�J�t�8 t@��I��u�8 ^u+D$Ë�ËT$V�t$3��2;�r;�sjX�T$^�
�V�t$W�|$V�7�6���������t�FPj�0��������t�F�FP�w�0��������t�F�FP�w�0������_^ËD$VW�0�x����0�4?���H�׉p�����_�H^ËD$VW�P�H�������ΉH��������_�P�^�U����ES�]3�;�V�E�N@  ��S�SvQW�E��}�S��p���S�j����E�PS����S�Z����E�e� �e� � �E��E�PS��������E�Mu�3�_9Su(�K�����C�����������E���  �s��Ӿ �  �suS������E���  Y��f�E�^f�C
[��U���\SVW�}�E�j�E�3�Z�E؉U�E��E��E܉E��EԉEЉE�E��E�}��� t��	t
��
t��uG��j^�G���w  �$� ��1|��9j�  :DBuj�F  �Ã�+tHHt����  �   j�E� �  X맃e� jX란�1�U�|��9~�:DB��   ��+t1��-t,��0tR��C��  ��E~��c�{  ��e�r  j��  Oj��  ��1|	��9�V���:DB�Y�����0��  �������U�9@B~��VP����YYjZ��LB�ÊA#ƅ�t�}�s�E��E���0�E���E��G�:DBug��������}� �U��U�u��0u�M��G��9@B~��VP����YYjZ��LB�ÊA#ƅ�t�}�s�E��E���0�E��M���G빀�+�
�����-���������9@B�U�~��VP诿��YYjZ��LB�ÊA#ƅ���   ���W�O���1�M|��9~D�Ã�+ttHHtd���  j�e�U���0u�G����1��   ��9��   �
��1|��9	j	XO������0uD���}  t*�ÍO���+�MtHH��   �M��jX����jX����j
OX��
��   �o����}�   �E�   3��=@B~��jP�þ��YY��LB�ÊA����t�ˍ��tAЁ�P  �G뾾Q  �u�=@B~��jP�y���YY��LB�ÊA����t�G��O����E�}� �8��   jX9E�v�}�|�E��E��E�H�E���E�}� ��   H�8 u�M��E���E�P�E��u�P�j����E�3Ƀ�9M�}��E�9M�uE9M�u+E=P  ~0�E�   �]�u�E�U�}� t`3۸�  �   �3��E�   �^=����}	�E�   ���uP�E�P��  �U��]uƋEʃ��3�3�3�3��3�3�3�3��E�   ��}� t3�3�3�3��E�   �ME�_�q�Yf�A
�E�^f�[�����q�����m�������Q�;��U����ES�]V�Ⱦ�  �� �  #�f��W�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   ��t�C-��C �}f��u��u9}uf�# �C �C�C0��  f;�uz�   �f� ;�u�} t��   @uh8)�Ff��t��   �u�} u.h0)�;�u#�} uh()�CP�H���Y�CY�e� �n  h )�CP�+���Y�CY���ϋ���i�M  ��f�e� j�Nf�U�k�M�}�����E���E�����P�E�P��
  ��f�}��?r�E�FP�E�P�  YY�Ef�3t�}�����������}��~j_�u����?  f�e� �E   �E�P�]����MYu��}�ށ��   ~�E�P�n���NYu�O�C�ɉE~P�M�u��}���E�P������E�P�����EP�E�P�����E�P������E��M�e� ��0�E�M�u��E�H�HH��5�K|0;�r�89u� 0H��;�s@f�� *�,�C���d �E�_^[��;�r�80uH��;�s�f�# �C �C�0�c jX�ӋL$V;��WsX�����<��������4������@t7�8�t2�=�}u3�+�tItIuPj��Pj��Pj��� ��0�3���(���� 	   �&����  ���_^ËD$;��s�ȃ����������D���t� ������� 	   ������  ���ËD$S�ȃ���VW�4��������<�����~ u#j�S����~ Yu�FP�� �Fj����Y��D8P�� _^[ËD$�ȃ����������D�P�� �SWj3������Yj_9=��~]V�h��������tA�@�tP�  ���YtC��|)�h���� P�H �h��4�����h�Y�$ G;=��|�^j�����Y��_[�V�t$V�#   ��Yt���^��F@t�v�  ��Y^��3�^�SV�t$3�W�F�ȃ���u7f�t1�F�>+���~&WP�v�������;�u�F��t$��F��N ����F�f �_��^[�j�   Y�SVWj3�3������3�Y95��~t�h�����t_�@�tYPV������h�YY���H���t0�|$uP�������YtC��|$ u��tP�������Yu��h��4�V�����YYF;5��|�j�����|$Y��t��_^[�V�t$;5��s@�΋������������D�t%WV�����t$�t$V�(   V�����������_^��G���� 	   �E����  ���^�U����e� �} S�]VW����  �E�ȃ����4������<�����ƊH����  ��Ht�@<
t�M���S�E�   �D0
�E�j P��uR�40�� ��u9�( j^;�u����� 	   �����0���m�$  P����Y����  ��U�U��L0�D0����   ��t	�;
u�$���E�M��E�;��M���   �E� <��   <t�C�E�   I9Ms�E@�8
u�E�^�C�E�s�E�j P�E�E�jP��40�� ��u
�( ��uG�}� tA��D0Ht�E�<
t��C�D1�);]u�}�
u�
�jj��u�������}�
t�C�M�9M�G������t0��@u�+]�]��E��3�_^[��S3�9�u�D$��a|Y��zT�� [�V��WV�� 9��=� tV��j�����Yj[�t$�   ��Y�D$t
j����Y�V�׋D$_^[�U��Q�=� Su�E��a��   ��z��   �� �   �]��   }(�=@B~jS�~���YY��LB�X����u���k�LB�������DJ�t�e
 �E�]	j�	�e	 �]jX�M�jj jQP�EPh   �5��[����� ��t���u�E���E��M����[���������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð���@Ë���   t�B:u�A
�t���   t�f���:u�
�t�:au�
�t����������������U��V3�PPPPPPPP�U�I �
�tB�$��u����A�
�tF�$s���� ^����U��V3�PPPPPPPP�U�I �
�tB�$��u�
�t
F�$s�F��� ^��U���$S�]V�uf�K
3�W�E�E܉E��E�f�F
����  3�#�#ʁ� �  f=���U��  f�����  f������  f���?w3��:f������u�E�Vu3�9Fu9u�o  3�f;�u�E�Su9Cu9u�F�F��k  �E��E��E��E   �E���} ~IƍK�E��E�M�E�E��M�� �	���M����QP�1�|�������t�E�f� �E��m��M�uȃE��E��M�} ��E�  f�} ~%�E�u�E�P�����E��  Yf�} �f�} 9�E��  f�} }+�E��E���E�t�E�E�P����KYu�}� t�M�f�}� �w�E�%�� = � u5�}��u,�e� �}��u�e� f�}���u�Ef�E� ��f�E���E���EދEf=�sf�M��f��M��N�M�Nf�F
�f����f ��   ��� ���& �~_^[��U���S� m3Ƀ�`9Mtc}�E�`n�؉E��`9Mu�Ef�9MtAVW�E��T�}��;�t'�@f�<� ��4�r�}�����M��u�V�u�r���YY3�9Mu�_^[��V�t$W����F@t�f �V�޿��V�   V���"�������_^�V�t$W����F�t4V����V���}  �v�  ����}�����F��tP�,����f Y�f ��_^�S�\$;��VWsr�����<����Ã��4�����D0tRS������Y�D0t)S����YP�� ��u
�( ���3���t�����0����� 	   ���S����Y����o���� 	   ���_^[�����������U��WVS�u�}���x u;����
�t.�F�'G8�t�,A<ɀ� �A��,A<ɀ� �A8�t������x����=� j ����j�����$   ��   3ې
�t'�F�G8�t�PS�|����؃��r�����8�t�������X�u	����
j��������[^_��U��WVS�M���   �u�}���x uN�A�Z� �I �&
�t!
�tFG8�r8�w�8�r8�w�8�uIu�3�8���   �������   ���   ����=� j ������j�����$   ��3�3ۋ����t#�tFGQPS苮���؃�聮����Y;�u	Iu�3�;�t	�����r��X�u	������j�������ˋ�[^_��V�t$;5��s8�΋������������D�tWV����V�(   V�����������_^��=���� 	   �;����  ���^�V�t$WV�
������Yt<��t��uj�����j�������Y;�YtV�����YP�� ��u
�( ���3�V�A����ƃ���Y�������d� ��tW�?���Y����3�_^�V�t$�F��t�t�v����f�f��3�Y��F�F^��%�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �+ �+ �+ �+ �+ , , *, 4, D, R, b, p, �, �, �, �, �, �, �, - "- <- R- j- �- �- �- �- �- �- �- �- . . . (. @. X. j. �. �. �. �. �. �. �. �. / / ,/ >/ N/ ^/ n/ z/ �/               �?    � 0 � 0N op O @N� �N�  N N o�mP;�m0N@N@Q�  O �O 0N o�S O @N� �N      �?   <  �@  �>          `@  �B         @�@      Y@:�0�yE>����Mb ?  @� P� Pf`f@N  �P� Pf`f@N�  !�!0N o�%O @N� �N  @+@N�m0N�)�m�m�m�m�m�m�m�m�m�n o o  @+@N�m0Np+�m�m�m�m�m�m�m�m�m�n o o  �,@N�m0N-�m�m�m�m�m�m�m�m�m�n o o@J N N0N o0NO @N� �H        pN N N0N o0NO @N� �N�O N N o�mQ�m0N@N@Q   k m@l m       �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    e+000          EEE50 P     (8PX 700WP        `h````  ppxxxx          ( n u l l )     (null)  __GLOBAL_HEAP_SELECTED  __MSVCRT_HEAP_SELECT    runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
abnormal program termination
    R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Microsoft Visual C++ Runtime Library    

  Runtime Error!

Program:    ... <program name unknown>  _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   modf    fabs    floor   ceil    tan cos sin sqrt    atan2   atan    acos    asin    tanh    cosh    sinh    log10   log pow exp ����    (�����    x�����    ;�����    ������    g�����    é�������             ��      �@      �        ����    ������    V�����    ������    C�GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll              ����!�%�    ������������5�9�1#QNAN  1#INF   1#IND   1#SNAN  H:mm:ss dddd, MMMM dd, yyyy M/d/yy  PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    �*         �/                        �+ �+ �+ �+ �+ , , *, 4, D, R, b, p, �, �, �, �, �, �, �, - "- <- R- j- �- �- �- �- �- �- �- �- . . . (. @. X. j. �. �. �. �. �. �. �. �. / / ,/ >/ N/ ^/ n/ z/ �/     � GetCommandLineA tGetVersion  >GetProcAddress  &GetModuleHandleA  � GetCurrentThreadId  �TlsSetValue �TlsAlloc  �TlsFree qSetLastError  �TlsGetValue GetLastError  } ExitProcess �TerminateProcess  � GetCurrentProcess mSetHandleCount  RGetStdHandle  GetFileType PGetStartupInfoA U DeleteCriticalSection $GetModuleFileNameA  � FreeEnvironmentStringsA � FreeEnvironmentStringsW �WideCharToMultiByte GetEnvironmentStrings GetEnvironmentStringsW  	GetEnvironmentVariableA uGetVersionExA �HeapDestroy �HeapCreate  �VirtualFree �HeapFree  �WriteFile RaiseException  �HeapReAlloc �HeapAlloc �HeapSize  �InterlockedDecrement  �InterlockedIncrement  jSetFilePointer  f EnterCriticalSection  �LeaveCriticalSection  �MultiByteToWideChar �InitializeCriticalSection � GetCPInfo � GetACP  1GetOEMCP  �VirtualAlloc  �LoadLibraryA  /RtlUnwind SGetStringTypeA  VGetStringTypeW  �LCMapStringA  �LCMapStringW  |SetStdHandle  ReadFile  � FlushFileBuffers   CloseHandle KERNEL32.dll            �LH    �/          �/ �/ �/ �q �/   Riptide.cdl c4d_main              �\�j        �w#�B�        ��                    riptide.tif redilogo.tif    At least one mesh object contains Ngons with 'holes'...

Click Yes to disable exporting Ngons and Continue.
Click No to Cancel. GetNgon() failed    InitObject() failed Riptide does not support "Shader" materials - using default.    Mem: m_pRegions[i].pFaceIndices _Rgn    Mem: m_pGroups[i].pFaceIndices  Mem: m_pRegions _Grp    Mem: m_pMats[i].pFaceIndices    Mem: m_pGroups  Mem: m_pMats    Mem: pRegionPolyCount   Mem: rgn_pPolymask  Mem: pGroupPolyCount    Mem: grp_pPolymask  Mem: pMatPolyCount  no NgonData Riptide Error: GetAndBuildNgon() failed #  http://skinprops.com
    #  Red-i Productions
   #  
    #  (a free plugin for Cinema 4D PC & Mac, R7.3 or later)
   #  Exported by Red-i Productions' "Riptide"
    #  Wavefront Material file
 #  ==========================================================================
  mtllib %s
  mtl disp %s
    map_d %s
   bump %s
    map_Ks %s
  map_Kd %s
  map_Ka %s
  Ks %f %f %f
    Kd %f %f %f
    Ka %f %f %f
    illum 2
    Ni %f
  d %f
   Ns %f
  newmtl %s
  
   Updating .mtl file...   newmtl %s   bump    map_d   map_Ka  map_Ks  map_bump    map_Bump    map_Kd  Ka %f %f %f Kd %f %f %f Ks %f %f %f Ni %f   Ns %f   disp     	  d %f    Setting up Materials... Riptide: Error parsing Ngon edges   Setting up Normals...   Setting up Group Tag... Setting up Region Tag...    Setting up Texture Coordinates...   Creating Polygon Object...  Polygon Object Allocation Failed    Creating Polygon Objects... default_Mat  %ld     %ld//%ld    %ld/%ld     %ld/%ld/%ld    f   f %ld %ld %ld %ld
  f %ld//%ld %ld//%ld %ld//%ld %ld//%ld
  f %ld/%ld %ld/%ld %ld/%ld %ld/%ld
  f %ld/%ld/%ld %ld/%ld/%ld %ld/%ld/%ld %ld/%ld/%ld
  f %ld %ld %ld
  f %ld//%ld %ld//%ld %ld//%ld
   f %ld/%ld %ld/%ld %ld/%ld
  f %ld/%ld/%ld %ld/%ld/%ld %ld/%ld/%ld
  # %ld facets

  usemtl %s
  # r %s
 g %s
   g %s %s
    Sorting by Material...  Sorting by Group... Sorting by Region...    Sorting by C4D Ordering...  # %ld texture coordinates

 vt %.08f %.08f
 BakeUVs failed  no uvTag    no UV Table no Texture Vertices # %ld vertex normals

  vn %.08f %.08f %.08f
   no Normal Vertex Table  no Normal Vertices  Ooops! Object named: %s has %d vertices, but zero faces!
No faces will be written.  Building tables...  no Faces    # %ld vertices

    v %.08f %.08f %.08f
    # r     g   %s %s   Processing:     #     (a free plugin for Cinema 4D PC & Mac, R7.3 or later)
    #  Wavefront OBJ format exported by Red-i Productions' "Riptide"
   Scanning Mesh...    obj Export .obj File    export.tif  %ld/%ld/     %ld/%ld/ %ld/%ld/ %ld/%ld/  %ld// %ld// %ld//  %ld  %ld %ld %ld    %ld/%ld  %ld/%ld %ld/%ld %ld/%ld    %ld/%ld/%ld  %ld/%ld/%ld %ld/%ld/%ld %ld/%ld/%ld    %ld//%ld     %ld//%ld %ld//%ld %ld//%ld default_Rgn default_Grp s %ld   usemtl %s   g %s    v %f %f %f  vn %f %f %f vt %f %f    mtllib %s   r %s    no Materials    no Regions  no Groups   no Vertices no Normals  no UVs  %ld/     %ld/ %ld/ %ld/ %ld//   no Index Data   no Segment Data Loading Mesh... Allocating Buffers...   Read Failed Scanning File...    Open Failed c4d Load Failed This plugin will only import Wavefront '.obj'
or '.mtl' format files - operation canceled.  OBJ MTL Import .obj File    import.tif  GroupTag.tif    RegionTag.tif   Txpmask dontXP.tif  res Riptide v1.9 .Obj Import/Export Plugin for C4D version R9.1 or later Installed. ==============================================================================      NOTREGISTRD Memory Allocation Error!
   Riptide: Memory Allocation Error -  File Error!
    Riptide: File Error -   u�  s�  �r�r�r    ��?          fmod         $x����t���������׭�������������������,$$ 	-]   ]       ����    ���� 
                                    �&   �&	   p&
   L&    &   �%   �%   �%   h%   @%   %   �$   �$x   �$y   �$z   x$�   t$�   d$   (    (   �'   �'   �'   �'!   �'   �'   �'   �'   �'   �'   �'   �'    �'   �'   �'   �'   �'   �'   x'   p'   h'   `'"   \'#   X'$   T'      �      ���������              �       �D        � 0                 ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ���d�j�o�u�z�������������ɯί�����>�C�]�b�������°����&�:�R�f���������ʱޱ��
�*�/�I�N�n�������βӲ���&�>�R�r�w�������ʳ�     .      VBVB                    ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                ���5      @   �  �   ����                     ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             H            `            0                                                                                                                          �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
       �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    PIPIhIhI���������   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   PI�                                   	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �           �&   �            C   C                                                                                                                                   C                                                                                                                                   l    `*\*X*T*P*L*H*@*8*0*$**** *�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)x)l)h)d)\)H)@)    .       �lH�H�H�H�H�H�H�H�H��l                     �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
�p     ����PST                                                             PDT                                                             �op����            ����        ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 0   000�01M1�1"2/2=2J2r2$3C4V4[4c4m4�;�;      L   d5h5l5p5t5x5|5�5�5�5�5�5�8�8�9�91:\:�:5;P;�;�;�;�;�<�<�=�=�=�>?�?�? 0  X   �0�01!2;2�2�2X3r354~4�4�45Q5s5�5�5H6j6�67r7�7
838u8�8�:T<x<�<p=�=�=D>�>,?U?�? @  H   *0s041e1�182m2�2�2%5^5�8�8�8t9�:�:�:>;k;�;E<�>�>�>�>�>�>�>�>�>   P  8   �3�3L9P9T9X9\9`9d9h9�<�=�=�=�=">L>v>�>�>�>c?�?   `  �   010?0Y0i0t0�0�0�0-1e1�1�1�1�1"2I2�2�2�23373c3�4�6�6�6�6�6�67�7�7�7�7�7�7�7@8E8\88�8�8�8�8�89$9J9O9t9y9�9�9�9�9!:o:�:;y;�;�;�;�;V<x<|<�<�<�<�<�<�< p  �   90�0�01:1X1v1�1�1�1�1
2,2J2h2�2�2�2�2�2)3G3e3�3�3�3�3�3444R4t4�4�4�4�4	5&5D5b55�5�5~6�6U7a7r7�7�7Q8�89�9@:�:;";:;l;�;�;�<�<�<b=�=�=�=�=�=�>�>�>?I?Y?i?z?   �  X   L0^0u01#1�1�11283�3F4�4�455@5)6[6�6�6�6R789�9*<�<�<�<=E=�=�=�=>0>M>a>?S?~? �  @   0o5�566a6F7�7	8�899:�:C;Z;u;�;�;S<_<p<�<�<�<�<�=�=>�> �  <   �3r4�4�4�56�67�7�859�9�9:!:e:#;-;>;`;�;�;�;r<�<8= �  8   �283�3�3�4�454667�7�8�9�<	=Z=�=3>�>�>_?�?�?   �  x   "0<0@0D0H0L0P0T0X0y0�1*2�2n3�344444 4$4(4I4K5�56�6$7H7L7P7T7X7\7`7d7�7J899�9:�:�:$;�;�<�<:=�=1>�>�>�?   �  �   C0Z0�0>1�1%2b23�3�3Q4�4H5�5?7]7u7�7�7�7!8�8�8�8�809>9L9]9�9�9�9:A:W:�:�:=;T;�;�;�;<�<�<�<�<==�=&>`>�>�>?)?J?�?�?�?�?�? �  �   000L0^0}0�0�0�0�0�01*1L1a1y1�1�1�1�112G2]2�2�2�2�233R3h3~34.4E4�4�4�45545�5�5�5�56-6T6k6�6G7�7�78*8S8p8�8�8@9o9�9�9�9&:@:�:A;q;�;�;�;�<�=r? �  l   l0�0-1\1�122�23L3�3a4�4�4�45B5l5�5�5�5�7�7�8�8�8=U=i=p=v=�=�=�=�=�=>>.>r>�>�>�>??S?X?�?�?�?   �   0020d0i0{0�0�0�0�0�0�01>1U1�1�1�1�1/2O2s2�2�2�2�23/3O3o3�3�3�3 44`4d4h4l4p4t4x4|45$5}5�5�5�5666Y6|6�67=7�7�7F8r89G:�:�:\>�>�>�>�>�>
??(?-?C?�?�?�?  �    0$0s0x0�0�071<1R1�1�1�1"2-262�2�2�2�2�3�3�3�3�4�4�4�4b5{5�5�5=6T6p6�6�67)7@7�7�7�7�7X8�8�8�8�8�8�809j9�9�9�9):^:�:�:�;R<�<�=>�>�>�?�?�?     D   }0�023#3�5�5�9�9�9�9�9�9�:�:�:.;A;�;8<F<`<�<�<=x=�=�=�=i> 0 �   �05�5r8�8�8/9�:\;j;�;�;$<H<l<�<�<=,=;=G=U=Z=d=v=�=�=�=�=�=�=�=�=�=�=�=�=�=>	>>>> >%>*>/>4>9>>>C>I>O>U>Z>_>e>j>p>u>z>>�>�>�>�?�?   @ �   D0�0�0�01&1Q1a1�1�1�1�1=2}2�2B3�3�3�34!4A4a4q4�4�4�4�45�5�5�5�5q6�6�6717Q7q7�7�7�7�7!8g8::#:j:r:�:�:
;K;�;�<(=Q={=�=�=�=Z>�>�? P �   0010Q0q0�0�0�1!313Q3�3�3 4J4�4e6Q7q7�7�7�7�7�78-8Q8�89!9Q9q9�9�9�9�9::1:Q:q:�:�:�:;�;�;�;�;E<�<�<�<=1=`=�=�=�=�=>A>Q>q>�>�>�>�>�>?@?�? ` �   0�0�0�0�0$1m1�1�1�1�1212Q2q2�2�2�23!313A3Q3�3�3�34T4�4�45I5�5�5�5�5�56�6R8Z8b8j8r8z8�8�89s9/:g:u:�:�:�:�:�:�:;H;M;q;�;�;<<!<b<q<�<�<=1=Q=>
>>>>&>->4>;>B>I>P>W>^>>?   p �   1'111;1�1�12=2Q22�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2333�5�5�5�5�5�5�5�56
66.6<6D6J6�6�6�67%7A7P7[7b7}7�7�7�7�7�7�7�7�7888(8\8e8�8�8�8�8�8�8�8�89k9f:r:�;3=;=�=�=E>T>j>�? � X   T0^1�1�1�1R255"5&5*5.5256546L6�6�6�8�8�89"969�9�95:[:k;z<�<f=}=�=�=z>�>�>�>�? �   *0G0C1K1e1k1|1�1�1�1�1�1�1�1�1�122(2A2�2�2�2�2�2�2�2�23+323B3H3O3Y3r3z33�3�3�3�3	4414E4w4~4�4�4�4�45)5S5a5�5�5�5�5�5�5	6;6K6�6�6�6�6�6�6�6�697@7�7�7�8�8�89 9,9<9{9�9�9:9:{:�:�:�:;�;�;�;�;�; <<<<$<K<W<_<g<w<�<�<�<�<�<�<�<�<
==(=O=^=�=�=�=�=�=>%>,> � �   J0t1z1�1�1�1�1�1�1�1�1-2p2X3�3^4p4�4�4�4�4+5�5�5�5�5
6�677B7H7a7�7�7�7�7�7�7�8�8�899$929�9�9�9:Q:�:K;[;g;y;�;�;�< =�=>h>�>�>�>�>8?`?   � <   e6�7�78�8�8�89a:|:�:q;{;�;E=T=�=�=�=�=�=>S>e>x>�> � �   G2]2�5 666666E6k6�6�6�6�6�6�6�6�6�6�6�6�6 77j7u7�7�7�7�7�7�7�78$8(8,8084888<8@8�8�8�8�8�8�899�9�9�9�9T:�:A;Y;n;�; <<$<><L<Z<e<y<<�<�<�<�<�<�<�<	=,=6=?=[=~=�=�=�=�=�=>!>'>;?C?I?Q?�?�?�? � 4  000G0M0]0x0g1t1?2D2�2�2�2+313?3y33�3�3�3�3�3�3�3�3�3�3�3�3�3444J4e4u4{4�4�4�4Q5W5�5�5�5�5�5�5�56)686Y6_6�6�6�6�6�6�6�6�6�6�6�67)737>7H7R7X7�7�7�7�7�7�7�7B8H8f8w8�8�8�8�8�8�8	99'959D9U9�9�9�9�9�9�9�9�9:5:<:@:D:H:L:P:T:X:�:�:�:�:�:;%;@;G;L;P;T;q;�;�;�;�;�;�;�;�;�;�;:<@<D<H<L<�<�<�=�=�=�=   � �   Q0W0^0k0r0z0�0�0�0�0�2�2�233+313A3L3^3q3|3�3�3�3�3�3�3�3�3�3�3�3�354�4�6�6�6�6�6
777!7'7,727B7K7e7v7|7�7�7�;�;�;�;�;�;<<<<"<+<�<�<�<�<�<�<�<�<=="=1=i=v=�=�=q>w>�>G?T?c?�? � �   0j0a2j2p2|2�2�2�2�2�2�2�2�2�2�23&3n3�3�3>4X4a4	6.636O6b6i6{6�6�6�6�6�6�6E7W7w7|7�7�7�7�7�7�7�7�7828R8�8�8�8[9�9�;�;)<�<�<�<�<=*=o=�=\>t>�>�>   �   00
000000"0&0*0.0�0�01(1�2�2�23J3^3�3�3�3�3�344 4I4V4[4h4t4.555N5�5�5�5�5Q6X6�6�6p7z788%8+818r8�8�8�89r<�<j=z=�=�=>V>\>j>�>�>D?J?X?�?�?�?     j0t0�0�0   D  �0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x388(848@8L8�8�8�8�8�8 99999   0 �   00000(00>4>8>@>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @ �   0000$0,040<0D0L0T0\0d0>1B1F1J1N1R1V1Z1^1b1f1j1n1r1v1z1~1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122
222222"2&2*2.22262:2L2P2�4�4747D7T7P9T9X9\9   ` x   p9 <<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< p    H0L0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        