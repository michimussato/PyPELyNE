MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���F���������|�J���ߚI���ߚ_��������������ߚX���ߚN���ߚM���Rich���        PE  L ��M        � !	  �  �      D�     �                         �                              � N   t (                            ` \3  `�                            � @            �                           .text   ��     �                   `.rdata  >   �  @   �             @  @.data   �4                      @  �.reloc  �?   `  @   &             @  B                                                                                                                                                                                                                                                                                                                                                                                                        ��  ��u��' ��������������������������������U��E�� t��t3�]ù`8�3 �����]ø   ]����U��p8V��H�QV�ҡp8�H�U�AVR�Ѓ���^]� U��p8V��H�QV�ҡp8�U�H�E�IRj�PV�у���^]� ����������U��p8�H�U�I(��VWR�E�P�ыp8�u���B�HV�ыp8�B�HVW�ыp8�B�P�M�Q�҃�_��^��]���U��p8�E�H�U �E��VWR�UP�ERP�A$���U��$R�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�,_��^��]��������������U��p8�P�E���   ��VWP�EP�E�P�ҋu���p8�H�QV�ҡp8�H�QVW�ҡp8�H�A�U�R�Ѓ�_��^��]� ������������U��p8�P�E�RP��VP�E�P�ҋuP����X �M��Y ��^��]� �������̡p8�P@�B,Q�Ѓ����������������U��p8���   �R|]��������������U��VW���Z �~������4X �M�E�U�NR�ωF�X �M�uX _��^]� �������������3��������������̸�������������U��V��j����F    �F    �Z j ����Z �N�X ���7Z �Et	V��` ����^]� ̋A�QPjRj �A�Ij PQ�5} ����U���SVW��� � �N���貣 �p8�H�A�V(R�Ѓ��N8�5 �Nh�.W �N|�&W �p8�Q���   P�B�Ѓ����   �W ���   ��V ���   ��V ���   ��V ���   ��V ��  ��V ��  ��V ��,  �V ��@  ���V ��T  ���V ����^�p8�Q�B$h%� �Nh�Ћp8�Q�B$h>� �N|�Ћp8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�H���   P�A�U�R�Ћp8�Q�J�E�P�у� j �M��#V �U�R���   �dV �M��LV j �M��V �E�P���   �CV �M��+V j �M���U �M�Q��  �"V �M��
V j �M���U �U�R��  �V �M���U j �M��U �E�P��,  ��U �M���U 3�P�M쉆h  ��l  ��p  ��t  �eU �M�Q���   �U �M��U �   ��|  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ǆx      �p8�B�P$h�� ���ҡp8�P��x  �R0PhM'  ���ҡp8�P��|  �R0Ph#'  ���ҡp8�P���  �R0Ph!'  ���ҡp8�P���  �R0Ph '  ���ҡp8�P���  �R0Ph"'  ���ҡp8�P���  �R0Ph$'  ���ҡp8�P���  �R0Ph%'  ���ҡp8�P���  �R0PhF'  ���ҡp8�P���  PhG'  �R0���ҡp8�P���  �R0PhH'  ���ҡp8�P���  �R0PhI'  ���ҡp8�P���  �R0PhJ'  ���ҡp8�P���  �R0PhK'  ����h�� �)� ���˅�tP�S _��^[��]áp8�P��x  �R0PhM'  �ҡp8�P��|  �R0Ph#'  ���ҡp8�P���  �R0Ph!'  ���ҡp8�P���  �R0Ph '  ���ҡp8�P���  �R0Ph"'  ���ҡp8�P���  �R0Ph$'  ���ҡp8�P���  �R0Ph%'  ���ҡp8�P���  �R0PhF'  ���ҡp8�P���  �R0PhG'  ���ҡp8�P���  �R0PhH'  ���ҡp8�P���  �R0PhI'  ���ҡp8�P���  �R0PhJ'  ���ҡp8�P���  �R0PhK'  ����_��^[��]������������V��T  ����R ��@  �R ��,  �R ��  ��Q ��  ��Q ���   ��Q ���   ��Q ���   ��Q ���   ��Q ���   �Q �p8�H�A���   R�Ѓ��N|�Q �Nh�Q �N8�0 �p8�Q�J�F(P�у��N�͝ ��^��� �����U��]�g� �������U���   V����� ��u^��]�SW����� �E̡p8�H�A�U�R�Ћp8�Q�J3�Sj��E�hd�P�у��U�R��迥 �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃�S�E�PjSj?h'  ����� �p8�Q�J�E�P�у�jS���
� jjjj���� �p8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ�S�M�QSjj?h'  ���W� �p8�B�P�M�Q�҃�jj���� Sjjj���� �p8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у�S�U�RSjj?h'  ����� �p8�H�A�U�R�Ѓ�jj���&� Sjjj���� �p8�Q�E�P�J�ыp8�B�PSj��M�h��Q�҃�S�E�PSjj?h'  ���s� �p8�Q�J�E�P�у�jj���� SSSS���8� h   h  < j?h'  ���к �M��N �p8�B�P4jhrdrb�M��ҡp8�H�A�U�R�Ћp8�Q�JSj��E�hT�P�у��U�Rh   h  ( j�E�PhD h'  ���M� �F$�p8�Q�J�E�P�у�h@���\����, Ph<��M��, P��x���R�@ ��P�E�P�0 ��P�M�Q�0 ���M��%- ��x����- �M��- ��\����- �U�SR�]< ����t�N$S�E�P� �M���, �M���M ���B� �p8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃�S�E�PSjj9h'  ���� �p8�Q�J�E�P�у�jj����� SSjS���� �p8�B�P�M�Q�ҡp8�H�ASj��U�h4�R�Ѓ��M�QSSj9h'  ���/� �p8�B�P�M�Q�҃�jS��谶 �p8�H�A�U�R�Ћp8�Q�JSj��E�h,�P�у��U�RSSj9h'  ���η �p8�H�A�U�R�Ѓ�jS���P� �p8�Q�J�E�P�ыp8�B�PSj��M�h$�Q�҃��E�PSSj9h'  ���m� �p8�Q�J�E�P�у���豿 ��調 �p8�B�P�M�Q�ҡp8�HS�Aj��U�h��R�Ѓ�S�M�QjSj9h'  ���&� �p8�B�P�M�Q�҃�jj���f� Sjjj���� SSh�  j8h'  ��胸 ���� �p8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у�S�U�RSjj	h&'  ��蘾 �p8�H�A�U�R�Ѓ�jj
���پ jjj
j���Z� �p8�Q�J�E�P�ыp8�B�PSj��M�h�Q�҃��E�PSSj	h''  ���� �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ��M�QSSjh='  ���c� �p8�B�P�M�Q�҃������ �p8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у�S�U�RSjj9h('  ���s� �p8�H�A�U�R�Ѓ�jj��贽 Sjj
j���6� �p8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃��E�PSSj	h)'  ���� �p8�Q�J�E�P�у�SSh�   j9�*'  W���ȹ �p8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ��M�Qh+'  �U�R�Ή}�]�蠺 �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃��E�Ph,'  �M�Q�Ή}�]��F� �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у��U�Rh-'  �E�P�Ή}�]��� �p8�Q�J�E�P�ыp8�B�M��PQ�ҡp8�H�ASj��U�h��R�Ѓ��M�Qh.'  �U�R�Ή}�]�蒹 �p8�H�A�U�R�Ѓ���觻 �p8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃�S�E�PSjj9h8'  ���"� �p8�Q�J�E�P�у�jj���b� jjjj���� �p8�B�P�M�Q�ҡp8�H�ASj��U�hp�R�Ѓ��M�QSSj	h9'  ���A� �p8�B�P�M�Q�҃�SSj9h:'  ���L� �p8�H�A�U�R�Ћp8�Q�JSj��E�hl�P�у�S�U�RSSj	h;'  ��色 �p8�H�A�U�R�Ѓ�SSj9h<'  ���� ���^� ���W� ���P� ���I� �p8�Q�J�E�P�ыp8�B�PSj��M�hd�Q�҃��E�P��诿 �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�hP�R�Ѓ��M�Qh3'  ���?� �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�h8�P�у��U�Rh4'  ���� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h �Q�҃��E�PhE'  ��蟿 �p8�Q�J�E�P�у����S� �p8�B�P�M�Q�ҡp8�H�ASj��U�h�R�Ѓ��M�Qh>'  ���E� �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у��U�Rh?'  ����� �p8�H�A�U�R�Ћp8�Q�E�P�J�ыp8�B�PSj��M�h��Q�҃��E�Ph@'  ��襾 �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ��M�QhA'  ���U� �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�hd�P�у��U�RhB'  ���� �p8�H�A�U�R�Ѓ���躽 �p8�Q�J�E�P�ыp8�B�PSj��M�hL�Q�҃��E�Ph5'  ��諽 �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h8�R�Ѓ��M�Qh6'  ���[� �p8�B�P�M�Q�҃����� �p8�H�A�U�R�Ћp8�Q�JSj��E�h �P�у��U�Rh7'  ���� �p8�H�U�R�A�Ѓ����F� �p8�Q�J�E�P�ыp8�B�PSj��M�h�Q�҃��E�P���̻ �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ��M�QhL'  ���\� �p8�B�P�M�Q�҃����� �p8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у��U�Rh#'  ���� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃��E�Ph!'  ��費 �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ��M�Qh '  ���b� �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у��U�Rh"'  ���� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃��E�Ph$'  ���º �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h��R�Ѓ��M�Qh%'  ���r� �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�h��P�у��U�RhF'  ���"� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h��Q�҃��E�PhG'  ���ҹ �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�hl�R�Ѓ��M�QhH'  ��肹 �p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�JSj��E�hP�P�у��U�RhI'  ���2� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h8�Q�҃��E�PhJ'  ���� �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h �R�Ѓ��M�QhK'  ��蒸 �p8�B�P�M�Q�҃����ַ �p8�H�A�U�R�Ћp8�Q�JSj��E�h�P�у��U�R���]� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h�Q�҃��E�PhC'  ���� �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�ASj��U�h �R�Ѓ��M�QhD'  ��蝷 �p8�B�P�M�Q�҃����� ���*� h'  V�N�<� �E�_[^��]���U���(S�   V��|  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ǆx      �Ja ���F  �p8�Q@WP�B,�Ћp8�Q�RP��h�� �M�Q����P�M��< �M���< �E썾@  P����< �M��< �p8�Q���   j hM'  ���Љ�x  �p8�Qj ;Ë��   h#'  �Q  ����PSh#'  ��茶 �p8�Q���   j h!'  ����PSh!'  ���d� �p8�Q���   j h '  ����PSh '  ���<� �p8�Q���   j h"'  ����PSh"'  ���� �p8�Q���   j h$'  ����PSh$'  ���� �p8�Q���   j h%'  ����PSh%'  ���ĵ �p8�Q���   j hF'  ����PShF'  ��蜵 �p8�Q���   j hG'  ����PShG'  ���t� �p8�Q���   j hH'  ����PShH'  ���L� �p8�Q���   j hI'  ����PShI'  ���$� �p8�Q���   j hJ'  ����PShJ'  ����� �p8�Q���   j hK'  ����PShK'  ���Դ �p8�Q���   j h#'  ���Љ�|  �p8�Q���   j h!'  ���Љ��  �p8�Q���   j h '  ���Љ��  �p8�Q���   j h"'  ���Љ��  �p8�Q���   j h$'  ���Љ��  �p8�Q���   j h%'  ���Љ��  �p8�Q���   j hF'  ���Љ��  �p8�Q���   j hG'  ���Љ��  �p8�Q���   j hH'  ���Љ��  �p8�Q���   j hI'  ���Љ��  �p8�Q���   j hJ'  ���Љ��  �p8�Q���   j hK'  ����_���  ^[��]Í�T  ���Љ�|  �p8�Q���   j h!'  ���Љ��  �p8�Q���   j h '  ���Љ��  �p8�Q���   j h"'  ���Љ��  �p8�Q���   j h$'  ���Љ��  �p8�Q���   j h%'  ���Љ��  �p8�Q���   j hF'  ���Љ��  �p8�Q���   j hG'  ���Љ��  �p8�Q���   j hH'  ���Љ��  �p8�Q���   j hI'  ���Љ��  �p8�Qj hJ'  �ϋ��   �Љ��  �p8�Q���   j hK'  ���Ћ�|  QSh#'  �Ή��  �ɱ ���  RSh!'  ��赱 ���  PSh '  ��衱 ���  QSh"'  ��荱 ���  RSh$'  ���y� ���  PSh%'  ���e� ���  QShF'  ���Q� ���  RShG'  ���=� ���  PShH'  ���)� ���  QShI'  ���� ���  RShJ'  ���� ���  PShK'  ���� _^[��]�������U���D�p8�P�B\SVW3��y|V3�V�ω]��Ѓ����   �I �p8�Q�RPV�E�P����P�M��B6 �M��Z6 j �M��6 �E�P�M���6 ��u P�M���5 �M�Q�M���e6 �E� ��t�E���t�MЃ���	6 ��t�M������5 �}� �M�u+F��5 �p8�B�P\j V���҃���N���_��^[��]���5 _��^[��]��������U���W���}���Y �E��u_��]�SV����E ���u��B �ءp8���   �Bj jS���Ћp8���   �B|�ǐ   W���Ћ��B �ˋ��B ������   ����   �	��$    ���p8�Q@�BW�Ѓ��u"�p8�A@�PV�E��҃��P�E��HV�у��p8�B@�HW�у��t"�p8�B@�E��@V�ЋM��Q��PV�҃��p8���   �B(���Ћ���t�p8���   �B(���Ћ����[����M��B �ˋ��B ������   ����   ���    �p8�Q@�BW�Ѓ��u"�p8�A@�PV�E��҃��P�E��HV�у��p8�B@�HW�у��t"�p8�B@�E��@V�ЋM��Q��PV�҃��p8���   �B(���Ћ���t�p8���   �B(���Ћ����[����u���!C Pj S���6C �p8�Q�M��BpSh�a  ���   �ЋM�Q����E ^[�   _��]���W�����   u�p8�P�Bpj hp ��  ��3�_�V�pW ����u^_Ë��[ �p8�QdVP�BX�Ћp8�Q����  ��tP�Bphp ��^�   _ËBpj hp ��^�   _����U���SV�E�WP����  �E��M��U��}��]�E��E�M��p8���U��Q�R4P�Ơ   h�a  ���ҡp8�P�B4Wh�a  ���Ћp8�Q�B4Sh�a  ���Ћp8�E��Q�R4Ph�a  ���ҡp8�P�E��R4Ph�a  ���ҡp8�P�E�R4Ph�a  ����_^�   [��]�������������U���8V�$V ����u�M��1 3�^��]� SW���DA ���p8���   �Bx���Ћp8�Q�J�؍E�P�ыp8�B�P�M�QS�ҡp8�P�RP��h�a  �E�P�M��P�M��D1 �M��\1 Wj(���2W j �M��1 �E�P�M��1 �Mȋ��21 ��t[�p8�Q�Blj Vh�a  �M��Ѕ�t>�p8���   j j �ȋBW�Ћp8���   �R|�E�P���ҋ��[@ P���SC �M���0 �p8�H�A�U�R�Ѓ��M�0 _[�   ^��]� �U����  SVW��3��uЉ}���T �؍M;�u�w0 _^3�[��]� �p8�P�RPh�a  �E�P��P�M��-0 �M��E0 W�M���/ �E�P�M��0 ��t��|  �E�t�E� �M��0 �}� ��   �p8�Q�B`W�M��Ѓ����   �p8�Q�RPW�E�P�M���P�M��/ �M���/ Sh0u  �M��y0 ����trVj(���U �p8�P���   j h1u  �M���P���  �p8�Q���   j h2u  �M���P����  �p8�Q���   j h3u  �M���P��� �M�G�8/ �p8�Q�B`W�M��Ѓ���/����p8�Q�RPh�a  �E�P�M��P�M���. �M���. �E�P�M���. �M���. j �M��. �M�Q�M��(/ �M���. ���  �p8�B�P`3�V�M��u��҃����  ��    �p8�P�RPV�E�P�M���P�M��R. �M��j. �p8�P�Blj Sh@�  �M��Ћ����x  �p8���   �B����=*� uE�MЃ��  u9Vj(����S �p8�B@�H,V�ыp8���B�P�����ҍE�P���I/ �p8���   �B����=� uE�MЃ��  u9Vj(���S �p8�B@�H,V�ыp8���B�P�����ҍE�P����. �p8���   �B����=× uE�MЃ��  u9Vj(���:S �p8�B@�H,V�ыp8���B�P�����ҍE�P���. �p8���   �B����=D� uE�MЃ��  u9Vj(����R �p8�B@�H,V�ыp8���B�P�����ҍE�P���,. �p8���   �B����=Dm uE�MЃ��  u9Vj(���|R �p8�B@�H,V�ыp8���B�P�����ҍE�P����- �p8���   �B����=�p uE�MЃ��  u9Vj(���R �p8�B@�H,V�ыp8���B�P�����ҍE�P���n- �p8���   �B����=�  u,�MЃ��  u Vj(���Q ShP�  �M���, P���� �p8���   �P����=  ��  �EЃ��  ��  Vj(���pQ �M��(+ �p8�Q@�J$�E�PV�ыp8�B�Pt��h`�  �M���h�  �� �������� �p8�QWP�B|�M��Ѝ� ������ �p8�Q�Btha�  �M���h�  ��H������� �p8�QWP�B|�M��Ѝ�H����� �p8�Q�Bthb�  �M���h�  ��8������N� �p8�QWP�B|�M��Ѝ�8����P� �p8�Q�Bthc�  �M���h�  ��(������� �p8�QWP�B|�M��Ѝ�(����
� �p8�Q�Bthd�  �M���h�  �M������ �p8�QWP�B|�M��ЍM���� �p8�Q�Bthf�  �M���h�  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Q�Bthk�  �M���h�  �M����?� �p8�QWP�B|�M��ЍM��D� �p8�Q�Bthl�  �M���h�  ����������� �p8�QWP�M�B|�Ѝ�������� �p8�Q�Bthm�  �M���h�  �M����� �p8�QWP�B|�M��ЍM��� �p8�Q�Bthn�  �M���h�  ���������v� �p8�QWP�B|�M��Ѝ������x� �p8�Q�Bth��  �M���h�  ��p������0� �p8�QWP�B|�M��Ѝ�p����2� �p8�Q�Bth��  �M���h  ��P�������� �p8�QWP�B|�M��Ѝ�P������ �p8�Q�Bth��  �M���h~  ��`������� �p8�QWP�B|�M��Ѝ�`����� �p8�Q�Bth��  �M���h�  ���������^� �p8�QWP�B|�M��Ѝ������`� �p8�Q�Bth��  �M���h�  ��P������� �p8�QWP�B|�M��Ѝ�P����� �p8�Q�Bth��  �M���h�  ��p�������� �p8�QWP�B|�M��Ѝ�p������ �p8�Q�Bth��  �M���h�  ��@������� �p8�QWP�B|�M��Ѝ�@����� �p8�Q�Bths�  �M���h�  ���������F� �p8�QWP�B|�M��Ѝ������H� �p8�Q�Btht�  �M���h�  ��0������ � �p8�QWP�B|�M��Ѝ�0����� �p8�Q�Bthu�  �M���h�  ��0������� �p8�QWP�B|�M��Ѝ�0����� �p8�Q�Bthv�  �M���h�  �� ������t� �p8�QWP�B|�M��Ѝ� ����v� �p8�Q�Bthw�  �M���h�  ���������.� �p8�QWP�B|�M��Ѝ������0� �p8�Q�Bthx�  �M���h�  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Q�Bthy�  �M���hp  ��`������� �p8�QWP�B|�M��Ѝ�`����� �p8�Q�Bthz�  �M���hq  �M����_� �p8�QWP�B|�M��ЍM��d� �p8�Q�Bth{�  �M���hr  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Q�Bth|�  �M���hs  ����������� �p8�QWP�B|�M��Ѝ�������� �p8�Q�Bth}�  �M���ht  ��@������� �p8�QWP�B|�M��Ѝ�@����� �p8�Q�Bth~�  �M���hu  �M����M� �p8�QWP�B|�M��ЍM��R� �p8�Q�Bth�  �M���hV  �M����� �p8�QWP�B|�M��ЍM��� �p8�Q�Bth��  �M���hW  �M������ �p8�QWP�B|�M��ЍM���� �p8�Q�Bth��  �M���hX  ��x������� �p8�QWP�B|�M��Ѝ�x����� �p8�Q�Bth��  �M���hY  ��h������D� �p8�QWP�B|�M��Ѝ�h����F� �p8�Q�Bth��  �M��Ћ�hZ  ��X������ �p8�QWP�B|�M��Ѝ�X���� � �p8�Q�Bth��  �M���h[  ��H������� �p8�QWP�B|�M��Ѝ�H����� �p8�Q�Bth��  �M���h`  ��8������r� �p8�QWP�B|�M��Ѝ�8����t� �p8�Q�Bth��  �M���ha  ��(������,� �p8�QWP�B|�M��Ѝ�(����.� �p8�Q�Bth��  �M���hb  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Q�Bth��  �M���hc  ��������� �p8�QWP�B|�M��Ѝ������ �p8�Q�Bth��  �M���hd  ���������Z� �p8�QWP�B|�M��Ѝ������\� �p8�Q�Bth��  �M���he  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Q�Bthe�  �M���hf  ����������� �p8�QWP�B|�M��Ѝ�������� �p8�Q�Bthg�  �M���hg  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Q�Bthh�  �M���hi  ���������B� �p8�QWP�B|�M��Ѝ������D� �p8�Q�Bthi�  �M���hh  ����������� �p8�QWP�B|�M��Ѝ�������� �p8�Q�Bthj�  �M���hv  ���������� �p8�QWP�B|�M��Ѝ������� �p8�Qhq�  �Bt�M���hw  ���������p� �p8�QWP�B|�M��Ѝ������r� �p8�Q�Bthr�  �M���hx  ��x������*� �p8�QWP�B|�M��Ѝ�x����,� �p8�Q�Bth��  �M���hk  ��h�������� �p8�QWP�B|�M��Ѝ�h������ �p8�Q�Bth��  �M���hj  ��X������� �p8�QWP�B|�M��Ѝ�X����� �p8�Q@�J(j�E�PV�у��M��� �u�F�M؉u��� �p8�B�P`V�M��҃�������M�� �M� _^�   [��]� ��������U���   S�A �؍M��u�c 3�[��]� �p8�P�RPVh�a  �E�P��P�M�� �M��2 j �M��� �E�P�M��| �M��� ���  �p8�Q�B`W3�W�MЉ}��Ѓ����  ���$    �p8�Q�RPW��|���P�M���P�M�� ��|���� �p8�P�Blj Sh�8 �M��Ћ��u���`  Vj(���dB jS��� ��   �}��p8�Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Q���   j h�8 �M��Ћp8�E��Qj h�8 �M싂�   �ЍM�Q�M�S�E�� jj ���� �p8���   �Pj j���ҋ}�G�M�}��" �p8�P�B`W�M��Ѓ���(���_�M��� �M�� ^�   [��]� ����������U���(V�? ���M��u�� 3�^��]� �p8�P�RPWh�a  �E�P��P�M��} �M�� j �M��K �E�P�M��� �M؋��u ��t/Vhp �M��# �΋��B �p8�Qdj WP��  �Ѓ��M��: �M�2 _�   ^��]� �����U���SW�}�م���  V�EjP��� �M��� �p8�Q��p  �R$P�M��ҡp8�P�BpWh�8 �M��Ћp8��Q�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F �R0Ph�8 �M��ҡp8�P��p  �RD�E�PQ���   ����p  �p8���   �B4���ЋMPQ�������p8���   �P(���ҍM��� ���s���^_[��]� ����U��V�u��� �Mj ��� �p8�QP�BphP�  ���Ћ�^]� �����������U���4SV�uW��� �M�� �p8�H@�]�A$�U�RS�Ћp83����E��E�QP���   h�  �M��Ћp8�E��   �}��Q���   �E�Ph`�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Pha�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q�E����   Phb�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phc�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phd�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phf�  ���ҡp8���   �U�R��Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phk�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phl�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phm�  ���ҡp8���   ��U�R����p8�QQ�$h�  �M̋��   ���]��p8�E�   �Q���   �E�Phn�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R����p8�Q���   Q�$h  �M����]��p8�E�   �Q���   �E�Ph��  ���ҡp8���   ��U�R����p8�Q���   Q�$h~  �M����]��p8�E�   �Q�E����   Ph��  ���ҡp8���   ��U�R����p8�Q���   Q�$h�  �M����]��p8�E�   �Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   �U��R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phs�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Pht�  ���ҡp8���   ��U�R�Ћp8�Q��j h�  �M̋��   �Ћp8�E��}��Q���   �E�Phu�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phv�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��}��Q���   �E�Phw�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h�  �M��Ћp8�E��E�P�}��Qhx�  ���   ���ҡp8���   ��U�R�Ћp8�Q���   ��j hp  �M��Ћp8�E��}��Q���   �E�Phy�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hq  �M��Ћp8�E��}��Q���   �E�Phz�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hr  �M��Ћp8�E��}��Q���   �E�Ph{�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hs  �M��Ћp8�E��}��Q���   �E�Ph|�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j ht  �M��Ћp8�E��}��Q���   �E�Ph}�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hu  �M��Ћp8�E��}��Q���   �E�Ph~�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hV  �M��Љ}��p8�E��Q���   �E�Ph�  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hW  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hX  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hY  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hZ  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h[  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j h`  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q�����   j ha  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hb  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hc  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j hd  �M��Ћp8�}��E��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ћp8�Q���   ��j he  �M��Ћp8�E��}��Q���   �E�Ph��  ���ҡp8���   ��U�R�Ѓ�j �M�Qhf  �M��� P���w �M��� he�  �M���� �p8�B�@|�M�Q�U�R���ЍM���� j �M�Qhg  �M��� P���' �M���� hg�  �M��� �p8�B�M�Q�U��@|R���ЍM��� j �M�Qhi  �M��o� P���� �M��� hh�  �M��R� �p8�B�@|�M�Q�U�R���ЍM��R� j �M�Qhh  �M��� P��� �M��/� hi�  �M��� �p8�B�@|�M�Q�U�R���ЍM��� j �M�Qhv  �M���� P���7 �M��߿ hj�  �M��� �p8�B�@|�M�Q�U�R���ЍM�貿 j �M�Qhw  �M��� P���� �M�菿 hq�  �M��b� �p8�B�@|�M�Q�U�R���ЍM��b� j �M�Qhx  �M��/� P��� �M��?� hr�  �M��� �p8�B�@|�M�Q�U�R���ЍM��� j �M�Qhk  �M���� P���G �M��� h��  �M���� �p8�B�@|�M�Q�U�R���ЍM��¾ j �M�Qhj  �M��� P���� �M�蟾 h��  �M��r� �p8�B�@|�M�Q�U�R���ЍM��r� �p8���   �
�E�P�у��M�� _��^[��]� ��������U��V�u���" �p8�H@�U�A$VR�Ѓ���^]� ������U���LSV��W�M��� �p8�H�A�U�R�Ѝ~�����OT �Mȋ��� 3�����   �M�Q�U�RV���KT �p8�P�Bth0'  �M��Ћp8���   P�B8�Ѓ�����   �p8�Q�Bth/'  �M��Ћp8���   P�BH�Ћp8�Q�R�M�QP��3��E�E��p8���   �I$�U�R�E�P�ыp8�B���   ���M�QV�M��ҡp8���   ��U�R�Ѓ�F;��'����p8�Q�B`j �M��Ћu�΃��u#j �� �M�� �p8�Q�J�E�P���"�U�R�� �M��� �p8�H�A�U�R�Ѓ��M��� _��^[��]� ����������U���xSVW�M��O �p8�H@�]�A$�U�RS�Ћp8�Q�B`��3�W�M��Ћ����t*V�M��� =�   tZ�p8�Q�B`GW�M��Ћ����u֋p8�Q�u�BV�Ћp8�Q�Bj j�h��V�Ѓ��M�� _��^[��]� �M���  �p8�Q���   PV�E�P�M���P�M���  �M����  �M����  �E�P�M���  �M�Q�M��?�  �p8�RP�B<V�M��ЍM���  �p8�Q@�J(j�E�PS�ыp8�B�u�HV�ыp8�B�P�M�VQ�ҡp8�H�A�U�R�Ѓ��M��N�  �M��F _��^[��]� �����������U���   W3��}��\( ;�u3�_��]Ëp8�Q@SP�B,�Ћp8�Q�RP��h%� ��t���Q����P�M�� ��t����� W�M�� �E�P�M��   �� ��u"W�M��g �M�Q�M��   �� �E� ��t�E���t�M؃���z ��t�M��m �}� t�M��_ [3�_��]�V�M��� �p8�B�P`W�M��}��}��҃���9  �p8�Q�RPP�E�P�M���P��t����� �M�� �p8�P�RPh�a  �E�P��t�����P�M�� �M��� j �M�� �E�P�M��  �M؋�� ���[  �p8�Q�B`3�V�M��u��Ѓ���;  �p8�Q�RPV��`���P�M���P�M��L ��`����a �& �p8�Qj P�Blh@�  �M��Ѕ���   �p8���   �ȋB��=�  ��   �X& �p8�Qj P�BlhP�  �M��Ћp8�Q3��؋B`W�Mĉ}��Ћ����tE�& �p8�Qj P�BlV�M���;�u�E�   �p8�Q�B`GW�M��Ћ����u��}� u�p8�Q�u�BpSV�M���F�u�u�F�M؉u��q �p8�Q�B`V�M��Ѓ��������}�G�M��}��G ��t����< �p8�Q�B`W�M��Ѓ���������t)�M��  �E�    �I% ���b �؅�u,�M���  �M���  �M���  ^[3�_��]��	��$    ���p8�Q�B`3�V�Mč~�Ѓ��t6�d$ ��$ PV�M�� ;�u3��p8�Q�B`FV�M��Ѓ��uӃ�u�p8�Q�u��BpSV�M���F�u��p8���   �B(���Ѕ�t�p8���   �B(���Ћ��c���3��3 �g$ ����% �p8�Q�B`V�M��Ѓ��tK�D$ PV�M���  Pj-�E��/$ ����% �}� t�M�Q�  ���p8�B�P`FV�M��҃��u���# ���r% j �3 ����# ��� �M���  �M���  �M���  ^[�   _��]���������U��Q�# �E���u��]� �p8�P�M�BTVh�a  �Ћ���u^��]� �p8�Q�B`SW3�W���Ѓ��t?�]�p8�QP�BT���ЋM�Qh0u  ����  ;�t"�p8�B�P`GW���҃��u�_[3�^��]� _[�   ^��]� �����U��Q��" �E���u��]� �p8�P�M�BTVh�a  �Ћ���u^��]� �p8�Q�B`SW3�W���Ѓ��tI�]�p8�QP�BT���Ћp8�Q�M��Rlj Qh@�  ����;�t!�p8�P�B`GW���Ѓ��u�_[3�^��]� _[�   ^��]� �����������U��Q�7" �E���u��]� �p8�P�M�BTVh�a  �Ћ���u^��]� �p8�Q�B`SW3�W���Ѓ��tI�]�p8�QP�BT���Ћp8�Q�M��Rlj Qh�8 ����;�t!�p8�P�B`GW���Ѓ��u�_[3�^��]� _[�   ^��]� �����������U���SV���q! ��u�uj �����  ��^[��]� ���P ����t�W�M���  �EVP��3�������u�p8�QVP�Bp�M��п   ��$    �p8���   �B4���Ѕ�t�p8���   �B4�<���    �p8���   �B(���Ћp8���   ��u�B0���Ћ���u��5�B(���ЋM��VQ���������u�p8�B�PpVW�M���G���j����u�E�P����  �M��$�  _��^[��]� ���������U���V�M��A  ��u�uP����  ��^��]� W���! ����u�uP����  _��^��]� S�M��]�  �ϻ   �E�    �
� ����tD�E�M�VP������؅�u�p8�Q�E��RpVP�M����E��p8���   �B(���Ћ���u��p8���   �B4���Ѕ�ty�p8���   �B4���Ћ����� ������   �MVQ�M��V����؅�u�p8�M��B�PpVQ�M����E��p8���   �B(���Ћ���u��   ���$    ��p8���   �B(���Ћp8���   �υ�u�B0�Ћ���u��`�B(�Ћ������ ����tD�MVQ�M������؅�u�p8�M��B�PpVQ�M����E��p8���   �B(���Ћ���u���������u�M�Q����  �M��(�  [_��^��]� �������������U���V�M��A ��u�uj ����  ��^��]� ���# ��t��p8���   �ȋBX�Ћ���t�SW�M��Z�  �]�M�VS3�������u�p8�QVP�Bp�M��п   �p8���   �B4���Ѕ�t�p8���   �B4�<��$    �p8���   �B(���Ћp8���   ��u�B0���Ћ���u��3�B(���ЋM���VS������u�p8�Q�BpVW�M���G���l����u�M�Q�����  �M����  _[��^��]� ����������U���V� ����u�uP���s�  ��^��]� �M��B�  ���k" ��u�uP���L�  �M���  ��^��]� �p8���   �ȋBXW3��Ћ���u�uP����  �M��L�  _��^��]� �p8�Q@�BV�Ѓ��t�p8�Q�BpVj �M��п   �I �p8���   �B4���Ѕ�t�p8���   �B4�=���    �p8���   �B(���Ћp8���   ��u�B0���Ћ���u��;�B(���Ћp8�Q@���BV�Ѓ��t�p8�Q�BpVW�M���G���c����u�M�Q���E�  �M��]�  _��^��]� ���j j j j�j�h%� j���J � ����U��EPj h%� ����o ]� ������U��p8�P�B`��\SVW��3��_hV���Ѓ����   ��|�}���p8�Q�M��RPV�E�P��P�M���  �M���  �p8�H�A�U�R�Ћp8�Q���   ���E�Ph N  �M�Q�M��ҋ��p8�H�A�U�R�Ћp8�Q�J�E�PW�ыp8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�Rx���EP�M��҅�tW�p8�H�A�U�RF�Ѓ��M���  �p8�Q�B`V���Ѓ�������p8�Q�J�EP�у�_^3�[��]� �p8�B�P�M�Q�҃��M���  �p8�H�A�UR�Ѓ�_^�   [��]� ���������U��p8�P�B`��XSVW�y|3�V���Ѓ���   ���$    �p8�Q�RPV�E�P����P�M���  �M��*�  �p8�H�A�U�R�Ћp8�Q���   ���E�Ph N  �M�Q�M��ҋءp8�H�A�U�R�Ћp8�Q�J�E�PS�ыp8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�Rx���EP�M��҅�tW�p8�H�A�U�RF�Ѓ��M��s�  �p8�Q�B`V���Ѓ���	����p8�Q�J�EP�у�_^3�[��]� �p8�B�P �M��ҋ�p8�H�A�U�R�Ѓ��M��
�  �p8�Q�J�EP�у�_��^[��]� ����������VW��� ����u_^Ë�Ǉp      � ��t�p8���   �ȋBX��PV���}���_�   ^������U���4SVW��� ' � ��� �p8�H�Q����W�ҡp8�H�A�UWR�Ѓ�����������~ ��u �p8�Q�J�EP�у�3�_^[��]� �p8�J@�Q,P�ҋp8�Q�RP��h%� �M�Q�ȉE���P�M����  �M����  �E��^hP�����  �M����  ���  u3�p8�Q�RP���e�W�E�P���ҋM�P�x�  �M���  �������p8�P�RP���e�W�E�P���ҋM�P�F�  �M��^�  ���������  u2�p8�P�RP���e�W�E�P���ҋM�P��  �M��#�  ���<������  u2�p8�P�RP���e�W�E�P���ҋM�P���  �M����  ���a����p8�P�M��BTh>� �E�    �Ћp8�Q�؋B`j �ˉ]��Ѓ����   ��I �]�p8�Q�E��R`P���ҋ��p8�P�BTW���Ћp8�Q���E��B��S�Ћp8�Q�J�ESP�у���������M�;�u�p8�B�P0jh�a  �����t�p8�P�B0j h�a  �ЋE��p8�Q�M�@�E�P�B`�Ѓ���K����& ��� j��$ �p8�Q�J�EP�у�_^�   [��]� �����U���(SV��MW��� �M���3�  �   ����  ��    �p8���   �B����=�  ��   9��  ��   �M����  j ���� �p8�QP�BphP�  �M��ЍM�Q�M��3�  �M���  ��t  �p8�RP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=  uy9��  uqW�M�Q���j���P�M���  �M���  ��t  �p8�RP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=*� ��   9��  ��   �M���  �p8�Q@�J$�E�PW�у��U�R�M����  �M����  �p8��t  �QP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=� ��   9��  ��   �M����  �p8�Q@�J$�E�PW�у��U�R�M��C�  �M��+�  �p8��t  �QP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=× ��   9��  ��   �M��F�  �p8�Q@�J$�E�PW�у��U�R�M���  �M��|�  �p8��t  �QP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=D� ��   9��  ��   �M���  �p8�Q@�J$�E�PW�у��U�R�M����  �M����  �p8��t  �QP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=Dm ��   9��  ��   �M����  �p8�Q@�J$�E�PW�у��U�R�M��6�  �M���  �p8��t  �QP�B$�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q��t  �RD�M�QP��,  ���t  �p8���   �B����=�p ��   9��  ��   �M��9�  �p8�Q@�J$�E�PW�у��U�R�M���  �M��o�  �p8�P��t  �R$P�M��ҡp8�P�BpWh@�  �M��Ћp8�Q��t  �RD�E�PQ��,  ���t  �p8���   �B(���Ћ���������M����  _^��[��]� ��������������U����   SVW�M�� ������  ����  �p8�Q@P�B,�Ћp8�Q�������   j h�  ���Ћp8�Qh�   �؋B4h�  ���Ћp8�Q���   j h�  ���Ћp8�Qjx�E܋B4h�  ���Ћp8�Q���   j h�  ���Ћp8�Qj�EЋB4h�  ���Ћp8�Q���   j h�  ������p8�]���EԍE��]�P�Q���   h�  ��D���Q���ҋ�M��P�U��H��M��P�]���p8�]��U���D����P���   �E�Ph�  Q���ҋ�M��P�UċH�MȋP�p8�ŰP�B4jh�  ���Ћp8�Q���   j h�  ���Ћp8�Qj �E�B0h�  ���Ћp8�Q���   j hR  ���Ћp8�Qj �E��B0hR  �����2� �E���u&�M�Q�2� ���E�    �M���  3�_^[��]� �p8���   �j h   ���ҋȉE����  �M����(�  �p8�H@�A$�U�RW�Ћp8�Q���   ��j h�  �M��Ћp8�Qj �����   h�  �M��ЋM�j jWP��� �}����U���R���  �E�WP��p����\���3�WW��p����M�  �M؁��   Q��8����h�  P�UR��T���P�7�  ����8������  �p8�Q�J�E�P�ыp8�BW�Pj��M�ht�Q�҃��E�P��T����;�  �p8�Q�J�E�P�ыM���jWhL  ��T���R�� �E�P���  �p8�Q�B4��Sh�  ���Ћp8�E܋Q�R4Ph�  ���ҡp8�P�EЋR4Ph�  ���ҡp8�P�EԋR4Ph�  ���ҡp8�P�R@�E�Ph�  ���ҡp8�P�R@�E�Ph�  ���ҡp8�P�E�PhR  �R0���ҡp8�P�E�R0Ph�  ���ҍ�T�����  j��p���ǅp�������|����}����  W��p�����  �M��U�  ��p����z�  �M��B�  �E�P�� ���M�}��+�  �G_^[��]� ���������������U��� SW�}�م���   V���$    ��p8�H�A�U�R�Ћp8�Q�Jj j��E�hx�P�у����� �p8�R�Rx�M�Q���ҋ�p8�H�A�ލU��RF�Ѓ���t!W�M�Q�������p8�B�P�M�Q�҃��p8���   �B4����P���<����p8���   �B(���Ћ����?���^_[��]� ������U���   SVW�Eċ�P�}������A	 �E܅��b  �p8�Q@P�B,�Ћp8�Q���ȋBTh%� �Ћ؉]����.  �p8�Q�B`j �M��E�    �Ћ�����}  ��	��$    ���]��p8�Q�J��d���P�ыp8�B���   ����d���QV��T���R�M��Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A��T���R�Ћp8�Q�J��d���P�ыp8�B�H����V�ыp8�B�P�M�VQ�҃����Q����p8�QP�BT���Ћ��u���  �p8�Q�BTh�a  ���Ћ؅���  V�M�Q���H����p8�B�P`j �M��E�    �҃���  ��I �M�QP�M���  ������   �p8�B�P`3�V���҃��t��p8�P�B`FV���Ѓ��u�M���  �p8�Q�B$V�M��Ћp8�Q�BpWh0u  �M��Ћ��� �p8�QP�B4h1u  �M��Ћ��$� �p8�QP�B4h2u  �M��Ћ��V� �p8�QP�B4h3u  �M��Ћp8�Q�RD�E�PV���ҍM��r�  �u�E��p8�Q@�E�P�B`�M��Ѓ��������}��p8�Q�BTh�a  ���Ћ؅��E  V�M�Q�������p8�B�P`j �M��E�    �҃���p  �p8�Q�M܋Rlj QP�M��ҋ����)  �p8�P�B`3�V���Ѓ��t�I �p8�Q�B`FV���Ѓ��u�p8���   �B����=�  un�M��'�  j ���� �p8�QP�BphP�  �M��Ћp8�Q�B$V�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q�RD�E�PV���ҍM��!�  �p8���   �B����=  uRW�M�Q�M�������p8�B�P$V�M��ҡp8�P�BpWh@�  �M��Ћp8�Q�RD�E�PV���ҍM���  �p8���   �B����=*� ��   �p8���   �B����=� th�p8���   �B����=× tN�p8���   �B����=D� t4�p8���   �B����=Dm t�p8���   �B����=�p uc�M���  �p8�Q@�J$�E�PW�ыp8�B�P$��V�M��ҡp8�P�BpWh@�  �M��Ћp8�Q�RD�E�PV���ҍM���  �u�E��p8�Q@�E�P�B`�M��Ѓ��������}��p8�Q�BTh�a  ���ЉE�����  V��t���Q���M����p8�B�P`j ��t����E�    �҃����  ��$    �p8�Q�M܋Rlj QP��t����ҋ؅��o  �p8�P�u��B`3�W���Ѓ��t��p8�Q�B`GW���Ѓ��u�M�jQ����� �M���b�  �p8�B�P$W�M��ҡp8�P�BpSh�8 �M��Ћp8��Q�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�FP�R0h�8 �M��ҡp8�P�F �R0Ph�8 �M��ҡp8�P�M��RD�E�PW�ҍM���  �E�p8�Q@�E�P�B`��t����Ѓ���G����}��u�F��t����u��b�  �M��Z�  �M��R�  �p8�Q�J�E�P�ыp8�B�P`��V�M��ҋ����������M���  �   _^[��]Ëp8�Q�J�E�P�у��M����  3�_^[��]ÍM����  �p8�B�P�M�Q�҃��M����  3�_^[��]ÍM���  �M���  �p8�H�A�U�R�Ѓ��M���  _^3�[��]����U���xSVW�E�P�M������  ���}���O  �p8�Q@�B,W�Ћp8�Q���ȋBTh%� �Ћ؉]����  �p8���   ���   ��jP�ωE����  �p8�Q�B`j �M��E�    �Ћ������  �p8�Q�J�E�P�ыp8�B���   ���M�QV�U�R�M��Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�H����V�ыp8�B�P�M�VQ�ҋM�������p8�QP�BT���Ѕ���  �p8�Q�ȋBTh�a  �Ћ�����  �p8���   �M����   �E�    �ЉE����  ��  ���$    ��p8���   �E��M����   P�ҋ����|  �p8�P�B`j ���E�    �Ћ؃��tH�p8�Q�BTS���ЋM�Qh0u  ����  ;��z  �E�p8�R@�E�P�B`���Ћ؃��u��p8�Q�B`3�S���Ѓ��t�p8�Q�B`CS���Ѓ��u�M���  �p8�Q�B$S�M��Ћp8�Q�BpVh0u  �M��Ћ��ݪ �p8�QP�B4h1u  �M��Ћ��� �p8�QP�B4h2u  �M��Ћ��A� �p8�QP�B4h3u  �M��Ћp8�Q�RD�E�PS���ҍM��]�  �E�@;E�E�������]�p8�u��H�A�U�FR�u��Ћp8�Q�B`��V�M��Ћ�����3����}�p8���   ���   �E�P�у������  �M����  �   _^[��]Ëp8�Q�BTS���Ћ΋��ϩ �p8�QP�B4h1u  ���Ћ��� �p8�QP�B4h2u  ���Ћ��5� �p8�QP�B4h3u  ���������p8�H�A�U�R�Ѓ��M��N�  3�_^[��]Ëp8�Q�J�E�P�у��M��(�  3�_^[��]Ëp8�B�P�M�Q�҃��M���  _^3�[��]����������U���   SVW�E�P�M��x�����  ���u̅�u�M����  3�_^[��]Ëp8�Q@�B,V�Ћp8�Q���ȋBTh%� �Ћ��}ȅ�t��p8���   ���   ��P�ΉE���  �p8���   �M䋂�   �Ћ؉]ą�t��p8�Q�B`j �M��E�    �Ћ������  ��I �p8�Q�J��|���P�у���|���RV�E�P�M��T}���p8�Q�J��|���P�ыp8�B�H����V�ыp8�B�P�M�VQ�ҋM܃��-����p8�QP�BT���Ћp8�Q�ȋBTh�a  �Ћ��u��E�    ����  �I �p8���   �E��M䋒�   P�ҋ��p8�P�B`j ���E�    �Ѓ���h  ���p8�QP�BT���Ћp8�Q�Rl�؋E�3�VPh@�  ����;��  ;���  �M���  �p8�P�B ���Ћp8�QP�B$�M��Ћp8���   �B����=�  ��   �M��B�  V���:� �p8�QP�BphP�  �M��ЍM�Q�M���  �M��o�  �p8�B�P`V�M�u��ҋ����tI�I �p8�P�BtV�M��Ћp8�QP���   V���ЋE��p8�Q@�E�P�B`�M��Ћ����u��p8���   �B����=  ��   W�M�Q�M�诼��P�M����  �M����  �p8�B�P`j �M��E�    �ҋ����tF�p8�P�BtV�M��Ћp8�QP���   V���ЋE��p8�Q@�E�P�B`�M��Ћ����u��p8���   �B����=*� ��   �p8���   �B����=� tl�p8���   �B����=× tR�p8���   �B����=D� t8�p8���   �B����=Dm t�p8���   �B����=�p ��  �M��[�  �p8�Q@�J$�E�PW�у��U�R�M���  �M���  �p8�P�B`j �M��E�    �Ћ�����t  �p8�Q�BtV�M��Ћp8�QP���   V���ЋE��p8�Q@�E�P�B`�M��Ћ����u��(  �p8�Q�]؋B`j ���Ѓ��t��$    �p8�Q�B`FV���Ѓ��u�p8���   �B����=�  un�M��g�  j ���^� �p8�QP�BphP�  �M��Ћp8�Q�B$V�M��Ћp8�Q�BpWh@�  �M��Ћp8�Q�RD�E�PV���ҍM��a�  �p8���   �B����=  uRW�M�Q�M������p8�B�P$V�M��ҡp8�P�BpWh@�  �M��Ћp8�Q�RD�E�PV���ҍM����  �p8���   �B����=*� ��   �p8���   �B����=� tk�p8���   �B����=× tQ�p8���   �B����=D� t7�p8���   �B����=Dm t�p8���   �B����=�p uf�]؍M����  �p8�Q@�J$�E�PW�ыp8�B�P$��V�M��ҡp8�P�BpWh@�  �M��Ћp8�Q�RD�E�PV���ҍM����  �Eԋp8�Q�u�@�E�P�B`���Ѓ��������]ċE�@;ÉE��K����}ȋp8�uЋQ�J�E�FP�u��ыp8�B�P`��V�M��ҋ�����_����p8���   ���   �U�R�Ѓ��M��]�  _^�   [��]��U���   SVW�E���P�]�������q�  ���}����  �p8�Q@�B,W�Ћp8�Q���ȋBTh%� �ЉEԅ���  �M�Q�������p8�B�P`j �M��E�    �ҋ�����w  ��]Сp8�H�A�U�R�Ћp8�Q���   ���E�PV��x���Q�M��ҋ�p8�H�A�U�R�Ћp8�Q�J�E�PV�ыp8�B�P��x���Q�ҡp8�H�A�U�R�Ћp8�Q�B����V�Ћp8�Q�J�E�VP�у��������p8�R�M�P�BT�Ѕ���  �p8�Q�ȋBTh�a  �Ћp8�Q�؋B`j �M��E�    �Ѓ���4  ���    �p8�Qj WP�Bl�M��ЉE����`  jW���� �p8�Q���B`j ���E�    �Ћ����tX�d$ �p8�Q�BTW���Ћp8�Q�M��Rlj Qh�8 ���ҋp8�Q��;E���  �E�@�E�P�B`�Ћ����u��p8�P�B`3�W���Ѓ��t��I �p8�Q�B`GW���Ѓ��u�M��q�  �p8�Q�B$W�M��Ћp8�E��Q�RpPh�8 �M��ҡp8�P��R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F�R0Ph�8 �M��ҡp8�P�F �R0Ph�8 �M��ҡp8�P�RD�E�PW���ҍM���  �E�p8�Q@�E�P�B`�M��Ћ}����������p8�u��Q�J�E�FP�u��ыp8�B�P`��V�M��ҋ������������D�  �M��<�  �M��4�  �   _^[��]ËBTW�Ћp8�Q�R0���Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F�R0Ph�8 ���ҡp8�P�F �R0Ph�8 ���������p8�H�A�U�R����p8�Q�J�E�P�у��M���  �M���  _^3�[��]���U���<SVW�E�P�M������&�  ������  �p8�Q@�B,V�Ћp8�Q���ȋBTh%� �ЉE�����  ����  �؅�u=Ph���M���o���M�Q�F] �p8�B�P�M�Q�҃��M��i�  3�_^[��]áp8���   �B����j =�  u��p8�P�B`�M�3��Ћ������   ���    �p8�Q�J�E�P�у��U�RV�E�P�M��Zp���p8�Q�J�E�P�ыp8�B�H����V�ыp8�B�P�M�VQ�ҋM����6����p8�Q�M�P�BT�Ѕ�tv�p8�Q�ȋBTh�a  �Ћp8��t|�QS�ȋBphp �Ћp8�Q�J�E�PG�ыp8�B�P`��W�M��ҋ���������M��6�  �   _^[��]áp8�H�A�U�R�Ѓ��M���  3�_^[��]ËQ�J�E�P�у��M����  _^3�[��]������U����  SVW���}��
�  ���2  �p8�Q@P�B,�Ћp8�Q�RP����h>� �E�P�Ήu���P�M��i�  �M���  �E��_|P����  �M��k�  ������Q��������p8�B���   j h#N  ���҅���  �p8�P�RPh%� �E�P����P�M����  �M���  �E���hP����  �M����  �p8�Q�B`j ���E�    �Ћ�����_  ���    �p8�Q�RPV�E�P����P��<�����  �M���  �p8�H�A�U�R�Ћp8�Q���   ���E�Ph N  ��d���Q��<����҉E��p8�H�A�U�R�Ћp8�Q�M��R�E�PQ�ҡp8�H�A��d���R�Ћp8�Q�J�E�P�ыp8�B�PP��h"N  �M�Q��<�����P���������  �M����  �M���  �p8�P�B$V�M���3��E��p8�E����   �R$�E�P�M�Q�ҡp8�P���   ���E�Ph N  �M��ҡp8���   ��U�R�Ћp8�Q�RD��������Ph"N  �M��ҡp8�P�RD�E�PV���ҡp8�u��P�B0jFh#N  �ˉu��Ћp83���t�����|������   �J0��t���SP�ыp8�B���   ����t���Q�M�h>� �ҡp8���   ���t���R�Ѓ��M����  ��������  �p8�Q�J�E�P�у���<�����  �p8�B�P`V���ҋ����������}��_��3��]�� �E���~V���� F;u�|�p8�P�B`3ۃ�|S�ω]��Ѓ���[  ��p8�Q�B`S���Ћp8�Q�RPP�E�P����P�M����  �M����  �p8�H�A�U�R�Ћp8�Q���   ���E�Ph N  ��d���Q�M��ҋ�p8�H�A�U�R�Ћp8�Q�J�E�PV�ыp8�B�P��d���Q�ҡp8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�P��(�EЋRxP�M��ҋ�p8�H�A�ލU��R���Ѓ���t�E�p8�Q�J�E�PC�у��M����  �p8�B�P`S���҃���������P����k�  �p8�P�B`3�S�ω]��Ѓ���v  �p8�Q�B`S���Ћp8�Q�RPP�E�P����P�M��^�  �M��v�  �p8�H�A�U�R�Ћp8�Q���   ���E�Ph N  ��d���Q�M��ҋ�p8�H�A�U�R�Ћp8�Q�J�E�PV�ыp8�B�P��d���Q�ҡp8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�P��(�EЋRxP�M��ҋ�p8�H�A�ލU��R���Ѓ���t �p8�Q�u��R8�E�PV��P�����F�u��p8�H�A�U�RC�Ѓ��M��Q�  �p8�Q�B`S���Ѓ��������E�H����  �E��E���I 3�9u���  ��I �p8�Q�J������P�ыp8�B���   ��������Q�~W��d���R��P����Ћp8�Q�J�؍����P�ыp8�B�P�����QS�ҡp8�H�A��d���R�Ћp8�Q�R\��������P������ҋءp8�H�A�����R�Ћp8�Q�J�����PS�ыp8�B�P������Q�ҡp8�H�A�U�R�Ћp8�Q���E�P������VQ��P������   �ҋءp8�H�A�U�R�Ћp8�Q�J�E�PS�ыp8�B�P������Q�ҡp8�P�R\��������P�M��ҋءp8�H�A�U�R�Ћp8�Q�J�E�PS�ыp8�B�P������Q�ҡp8�P�Rx�������P�M��ҋءp8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�����R�A�Ћp8�Q�J�����P�ыp8�B�P������Q�҃�����  �p8�H�A������R�Ћp8�Q���   ��������PV�����Q��P����ҋءp8�H�A�U�R�Ћp8�Q�J�E�PS�ыp8�B�P�����Q�ҡp8�H�A������R�Ћp8�Q�J������P�ыp8�B���   ��������QW������R��P����Ћp8�Q�J�؍�,���P�ыp8�B�P��,���QS�ҡp8�H�A������R�Ѓ��p8�Q�R8��,���PV��P����ҡp8�H�A��,���R�Ћp8�Q�J������P�ыp8�B�P8���M�QW��P����ҡp8�H�A�U�R�Ѓ���;u��0����   )E�)E�����3�9}��v  �d$ �M�踽  �p8�Q�J������P�ыp8�B���   ��������QW��<���R��P����Ћp8�Q�J��������P�ыp8�B�P������QV�ҡp8�H�A��<���R�Ћp8�Q�R8��������Ph/'  �M��ҡp8�H�A������R�Ћp8�Q�J������P�ыp8�B�P`��3�S�������ҋ������  �p8�H�A������R�Ћp8�Q���   ��������PV��l���Q�������ҋ�p8�H�A�� ���R�Ћp8�Q�J�� ���PV�ыp8�B�P��l���Q�ҡp8�H�A������R�Ћp8�Q�J������P�ыp8�B���   ��������QW������R��P����Ћp8�Q�J����@���P�ыp8�B�P��@���QV�ҡp8�H�A������R�Ѓ��p8�Q�Rx��@���P�� ����ҋ�p8�H�A�ލ�@����RF�Ћp8�Q�J������P�у���t�p8�B�P0jh0'  �M��ҡp8�H�A�� ���RC�Ћp8�Q�B`��S�������Ћ�����J����p8�Q�J��d���P�ыp8�B���   ����d���QW������R��P����Ћp8�Q�؋BV�Ћp8�Q�BVS�Ћp8�Q�J������P�ы]������r����p8���B�P��d���Q�ҡp8�P�RP��V�E�P�K|��P��<���藺  �M�诺  �p8�P���   j h�a  ��<����Ћp8�Q�J��uN������P�ыp8�B�Pj j�������h��Q�ҡp8�P�R8��������Ph1'  �M��ҍ������L������P�ыp8�B�Pj j�������h��Q�ҡp8�P�R8��������Ph1'  �M��ҍ������p8�H�AR�Ћp8�Q�RP��h"N  ������P��<�����P�M�荹  ������袹  �p8�P���   j h�a  �M��ЍM����~�  �p8�Q�RPh"N  ������P��<�����P�M��5�  �������J�  �p8�P���   j h�a  �M��ЍM��E��%�  �p8�Q�RPh"N  ������P��<�����P�M��ܸ  ��������  �p8�P���   j h�a  �M��ЍM�������ɸ  �p8�Qh"N  ������P��<����RP��P�M�耸  ������蕸  �p8�P���   j h�a  �M��ЍM����q�  �p8�Q�RPh"N  ������P��<�����P�M��(�  �������=�  �p8�P���   j h�a  �M��ЍM��E���  �p8�Q�J(��|���SP�ыp8�؋B�P�M�Q�ҡp8�H�A�U�RS�Ћp8�Q�J��|���P�ыp8�B�PH��jj �M��ҡp8�H�A(V��\���R�Ћp8�Q�J�؍E�P�ыp8�B�P�M�QS�ҡp8�H�A��\���R�Ѓ���
�J  �p8�Q�J��0���P�ыp8�B�Pj j���0���h��Q�ҡp8�H�A(������VR�Ћp8�Q�J��������P�ыp8�B�P������QV�ҡp8�H�A������R�Ћp8�Q�J������P�ыp8�B�@������Q��0���R�Ћp8�Q�B<��8�������Ћp8�Q�RLj�j�������QP�������ҡp8�H�I�U�R������P�ыp8�B�P������Q�ҡp8�H�A������R�Ћp8�Q�J��0���P�у��p8�u��B�P(�����VQ�ҋءp8�H�A�����R�Ћp8�Q�J�����PS�ыp8�B�P�����Q�҃���
�K  �p8�H�A������R�Ћp8�Q�Jj j�������h��P�ыp8�B�P(������VQ�ҋ�p8�H�A��p���R�Ћp8�Q�J��p���PV�ыp8�B�P������Q�ҡp8�H�A������R�Ћp8�Q�R������P������Q�ҡp8�P�B<��8�������Ћp8�Q�RLj�j���p���QP�������ҡp8�H�I�����R������P�ыp8�B�P������Q�ҡp8�H�A��p���R�Ћp8�Q�J������P�у��p8�u��B�P(��,���VQ�ҋءp8�H�A�����R�Ћp8�Q�J�����PS�ыp8�B�P��,���Q�҃���
�K  �p8�H�A�����R�Ћp8�Q�Jj j������h��P�ыp8�B�P(������VQ�ҋ�p8�H�A��P���R�Ћp8�Q�J��P���PV�ыp8�B�P������Q�ҡp8�H�A��$���R�Ћp8�Q�R��$���P�����Q�ҡp8�P�B<��8��$����Ћp8�Q�RLj�j���P���QP��$����ҡp8�H�I�����R��$���P�ыp8�B�P��$���Q�ҡp8�H�A��P���R�Ћp8�Q�J�����P�у��p8������B�P(��L���VQ�ҋءp8�H�A��,���R�Ћp8�Q�J��,���PS�ыp8�B�P��L���Q�҃���
�K  �p8�H�A������R�Ћp8�Q�Jj j�������h��P�ыp8�B�P(������VQ�ҋ�p8�H�A��`���R�Ћp8�Q�J��`���PV�ыp8�B�P������Q�ҡp8�H�A��t���R�Ћp8�Q�R��t���P������Q�ҡp8�P�B<��8��t����Ћp8�Q�RLj�j���`���QP��t����ҡp8�H�I��,���R��t���P�ыp8�B�P��t���Q�ҡp8�H�A��`���R�Ћp8�Q�J������P�у��p8�B�P������Q�ҡp8�H�Aj j�������h��R�Ћp8�Q�J������P�ыp8�B�Pj j�������h��Q�ҡp8�H�A������R�Ћp8�Q�Jj j�������h��P�ыp8�B�P�����Q�ҡp8�H�A��@j j������h��R�Ћp8�Q�J��d���P�ыp8�B�@��d���Q�����R�Ћp8�Q�B<����d����Ћp8�Q�RLj�j������QP��d����ҡp8�H�A��D���R�Ћp8�Q�R��D���P��d���Q�ҡp8�P�B<����D����Ћp8�Q�RLj�j���,���QP��D����ҡp8�H�A������R�Ћp8�Q�R������P��D���Q�ҡp8�P�B<���������Ћp8�Q�RLj�j�������QP�������ҡp8�H�A�����R�Ћp8�Q�����P�������RQ�ҡp8�P�B<��������Ћp8�Q�RLj�j��M�QP������ҡp8�H�A��4���R�Ћp8�Q�R��4���P�����Q�ҡp8�P�B<����4����Ћp8�Q�RLj�j�������QP��4����ҡp8�H�A��T���R�Ћp8�Q�R��T���P��4���Q�ҡp8�P�B<����T����Ћp8�Q�RLj�j��M�QP��T����ҡp8�H�A������R�Ћp8�Q�R������P��T���Q�ҡp8�P�B<���������Ћp8�Q�RLj�j�������QP�������ҡp8�H�A�U�R�Ћp8�Q�R�E�P������Q�ҡp8�P�B<���M��Ћp8�Q�RLj�j������QP�M��ҡp8�H�A������R�Ћp8�Q�J��T���P�ыp8�B�P��4���Q�ҡp8�H�A�����R�Ћp8�Q�J������P�ыp8�B�P��D���Q�ҡp8�H�A��d���R�Ћp8�Q�J�����P�ыp8�B�P������Q�ҡp8�H�A������R�Ћp8�Q�J������P�ыp8�B�P�M�Q�ҡp8�H�Aj j��U�h��R�Ћp8�Q�J��t�����@P�ыp8�B�@��t���Q�U�R�Ћp8�Q�B<����t����Ћp8�Q�RLj�j��M�QP��t����ҡp8�P�R8��t���Ph2'  �M��ҡp8�H�A��t���R�Ћp8�Q�J�E�P�ыM����U�RW��  �p8�H�A�U�RG�Ћp8�Q�J��,���P�ыp8�B�P�����Q�ҡp8�H�A�����R�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�҃���<���迪  �M�跪  ;}�������M��6�  ��P���蛪  ������萪  _^[��]����������U���V���"& ��u^��]�W3�Wj�E�P���E� '  �}��~J Wj�M�Q���E�!'  �}��fJ Wj�U�R���E�"'  �}��NJ Wj�E�P���E�#'  �}��6J Wj�M�Q���E�$'  �}��J Wj�U�R���E�%'  �}��J WW�E�P���E�='  �}���I h���h  �Wjh���h  �h,'  �M�Q���E�*'  �}��^  WW�U�R���E�9'  �}��I �E�:'  �}���WW���T$�E��$hgnlf��� �\$������\$�T$�$P�U ��WW���T$�M��$hgnlf��� �\$�E�<'  ����}��\$�T$�$Q��� ���|k���M�脨  �p8�B�P4htxt h1'  �M��ҡp8�P�B4hkhc h0'  �M��Ћp8�Q�B4htxt h/'  �M��Ћp8�Q�B4htxt h2'  �M��ЍM�Qj�N���  �������M��\�  �G_^��]����U���   SV���~� �E�����  ��W���H�  �M���辧  3���~�E�P�M�QV���H�  F;�|�U�R����  ���p8�H�&  �A�U�R�Ѓ��M�Q�M��U�R3�W�H� ���]  �E�;E��7  �p8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�H�U��I(R��x���P�ыp8���B�P�M�Q�ҡp8�H�A�U�RV�Ћp8�Q�J��x���P�ыp8�B�P�M�Q�ҡp8�H�I�U�R�E�P�ыp8�B�P<��8�M��ҋp8�Q�RLj�j��M�QP�M��ҡp8�P�B<�M��Ћp8�Qj��RLj��M�QP�M��ҡp8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�҃��E�P�M�Q�M�GW�� ��������M����  �E��U�RP���<�  �p8�Q�Bth/'  �M��Ћp8���   P�BH�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ѓ��M����  �p8�Q�J�E�P�у��M��إ  �U�R�� ��_��^[��]� �u�QV�ҡp8�H�Qj j�h��V�҃��M�薥  �E�P�ݫ ��_��^[��]� �p8�Q�u�BV�Ћp8�Q�Bj j�h��V�ЍM�Q蜫 ����^[��]� ���������������U���V�uW�����L  S�]��$    ��|  ��   �M�蛤  �p8�P��l  �R$P�M��ҡp8�P�BpVh0u  �M��Ћ���u �p8�QP�B4h1u  �M��Ћ��	v �p8�QP�B4h2u  �M��Ћ��;v �p8�QP�B4h3u  �M��Ћp8�Q��l  �RD�E�PQ��  �ҍM��M�  ��|   u.j �M����  �p8�P�RD�E�Ph�a  ���   �ҍM���  V���^�����l  �p8���   �B4����PS�������p8���   �B(���Ћ��������[_^��]� �������U���   �E�VP���  ����  �M�Q���  ���ƹ  �M���  �U�R�M��B�  �E�P�M�趄  �p8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�H�A�U�R�Ћp8�Q�R�E�P�M�Q�ҡp8�P�B<�� �M��Ћp8�Q�RLj�j��M�QP�M��ҡp8�H�A�U�R�Ѓ��M�Q��l����R�  ��l���R�E��uPV��  ����l���谁  �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�A�U�R�Ѓ��M��p�  �M��h�  ��^��]� ���������������U���8V�E��P�M�軀  P�M�Q���o����uPV腄  ���M���  �M���  �p8�B�P�M�Q�ҡp8�H�Aj j��U�ht�R�Ѓ��M�Q��舃  �p8�B�P�M�Q�ҡp8�H�A�UR�Ѓ���^��]� ���������U���  SVW��3ۉ}ĉ]����  ���u�;���  �E�P���ݶ  �M����  �p8���   �Sh   ���ЉE�;���  P�<�  �M�Q�S�  �����I����p8�B�PhS�M�]��҅��  �p8�P�E��RhP�M�ҋp8���   P�BH�Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A��8���R�Ћp8�Q�JSj���8���h��P�ыp8�B�Px��$��8���Q�M��ҋ�p8�H�A�ލ�8����R���Ѓ�;���
  �p8�Q�B����V�Ћp8�Q�J�E�VP�у���苬���X�v  �L�  ���U�  �p8�J@�Q,P�ҋ�p8�P���   ��Sh�  ���Ћp8�E�ǅ(���   ��0����Q���   ��(���Ph�  ���ҡp8���   ���(���R���E����������U��\$�G\�$蓾 �p8���������������   �J,P������P�ыp8�B���   ��������Qh�  ���ҡp8���   �������R���E���\$��t����G`�$�� �p8���������������   �J,P������P�ыp8�B���   ��������Qh�  ���ҡp8���   �������R�Ѓ��p8�Q�J��H���P�ыp8�B�PSj���H���h��Q�҃�������P�M��~  �p8�Q�J���� ���P�ыp8�B�P�� ���QV�ҡp8�P�B<���� ����Ћp8�Q�RLj�j���H���QP�� ����ҡp8�H�A��@���R�Ћp8�Q�R��@���P�� ���Q�ҡp8�P�B<����@����Ћp8�Q�RLj�j��M�QP��@����ҍ�@���P��`�����{  P�MQ��h���R��  ����`����`|  �p8�H�A��@���R�Ћp8�Q�J�� ���P�ыp8�B�P������Q�ҡp8�H�A��H���R�Ѝ�h���jQ�`�  ����u��h���R��  ��;���  ��  ���&�  ���?�  ���u�;��  ��u��p8���   �B����=�� ��  �������5�  �p8�Q@�J$������PV�ыp8�B���   ��Sh�  �������ҋ�p8�P���   Sh�  ��������S���������sz  ��u_;��D  �������+z  �p8�Q���   Ph�  ��`���P��������P�M��z  ��`�����z  �E�P�������~  ��   ����   ������Q���  ����  hh���`�����y  P������R�E�P��}  ����`����z  �M��}  �p8�Q�J������P�ыp8�B�PSj�������hd�Q�҃�������P�M���|  �p8�Q�J������P�эU�R�E�P��`���Q�o}  ��P�������0}  ��`�����y  �M���y  ��������y  S�M��y  �M��U�R��������}  ��t������SP��  ����u���2��E�t�e���M��y  ����  �M��|  �p8�Q�J�����P�ыp8�B�Pj j������h��Q�҃������P�M�� z  �p8�Q�J����P���P�ыp8�B�P��P���QV�ҡp8�P�B<����P����Ћp8�Q�RLj�j������QP��P����ҡp8�H�A��0���R�Ћp8�Q�R��0���P��P���Q�ҡp8�P�B<����0����Ћp8�Q�RLj�j��M�QP��0����ҍ�0���P�M���w  �p8�Q�J��0���P�ыp8�B�P��P���Q�ҡp8�H�A�����R�Ћp8�Q�J�����P�эU�R�EP��`���Q�d{  ��h\��������1w  P��`���R������P�={  ����������w  ������jQ�!�  ����u������R�·  ���E�P������Q������R��z  �p8�H�A������R�Ћp8�Q�Jj j�������hd�P�у� ������R��������y  �p8�H�A������R�Ѝ�����jQ苆  ����uP������R������P�φ  ���������w  ��������v  ��`�����v  �M���v  ��������v  �������͗  �u��}�3ۋp8���   �B(���ЉE�;�������M��/y  �p8�Q�J��|���P�ыp8�B�PSj���|���h��Q�҃���X���P�M��w  �p8�Q�J���� ���P�ыp8�B�P�� ���QV�ҡp8�P�B<���� ����Ћp8�Q�RLj�j���|���QP�� ����ҡp8�H�A�����R�Ћp8�Q�R�����P�� ���Q�ҡp8�P�B<��������Ћp8�Q�RLj�j��M�QP������ҍ����P�������u  P��h���Q������R��x  ���������au  �p8�H�A�����R�Ћp8�Q�J�� ���P�ыp8�B�P��X���Q�ҡp8�H�A��|���R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�hX�Q�҃�$�E�P�������w  �p8�Q�J�E�P�у�hBF ������SR��  P��  �����5  �������t  ��h����t  �p8�u��H�A�U�FR�u��Ћp8�Q�Bh��V�M�Ѕ��B����;  ShP���|����x:��Sh��M��j:����|���Q�U�R�E�P�����Q�_\  ��P��X���R�O\  P�' �p8�H�A��X���R�Ћp8�Q�J�����P�ыp8�B�P�M�Q�ҡp8�H�A��|���R�Ѓ� ��h����s  �p8�Q�J�E�P�у��M��s  �M�w�  �M�os  3�_^[��]�0 Sh���M��9���U�R�' �p8�H�A�U�R�Ѓ��������.s  ��h����#s  �p8�Q�J�E�P�у��u�U�R�b�  V��  ���M���r  �M��  �M��r  _^�   [��]�0 ���U���0  SVW��3ۉ}ԉ]����  ���u�;�t:�E�P����  �M��)u  �p8���   �Sh   ���ЉE�;�u#�M��rr  �M�j�  �M�br  3�_^[��]�0 P�Q�  �M�Q�h�  �����^����p8�B�PhS�M�]��҅��Y
  ��p8�P�E��RhP�M�ҋp8���   P�BH�Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A������R�Ћp8�Q�JSj�������h��P�ыp8�B�Px��$������Q�M��ҋ�p8�H�A�ލ������R���Ѓ�;��	  �p8�Q�B����V�Ћp8�Q�J�E�VP�у���蟞���X�v  �`�  ���i�  �p8�J@�Q,P�ҋ�p8�P���   ��Sh�  ���Ћp8�E�ǅt���   ��|����Q���   ��t���Ph�  ���ҡp8���   ���t���R���E����������U��\$�G\�$觰 �p8�������������   �J,P�����P�ыp8�B���   �������Qh�  ���ҡp8���   ������R���E���\$�������G`�$�/� �p8���������������   �J,P������P�ыp8�B���   ��������Qh�  ���ҡp8���   �������R�Ѓ���  ����  ����  ���u�;��1  ����$    �d$ �u��p8���   �B����=�� ��  ��������  �p8�Q@�J$������PV�ыp8�B���   ��Sh�  �������ҋ�p8�P���   Sh�  ��������S���������2n  ��um;��R  ��,�����m  �p8�Q���   Ph�  �����P��������P�M��mn  ������n  �E�P��������q  �M��n  ��,�����   ����   ��0���Q諳  ��蔥  hh�������m  P��0���R�E�P�q  ��������5n  �M��p  �p8�Q�J������P�ыp8�B�PSj�������hd�Q�҃�������P�M��p  �p8�Q�J������P�эU�R�E�P�����Q� q  ��P��������p  ������m  �M��m  ��0����m  S�M���l  �M��U�R�������wq  ��t������SP��|  ����u���2��E�t�e���M��Fm  ����  �M���o  �p8�Q�J������P�ыp8�B�Pj j�������h��Q�҃��� ���P�M��m  �p8�Q�J����l���P�ыp8�B�P��l���QV�ҡp8�P�B<����l����Ћp8�Q�RLj�j�������QP��l����ҡp8�H�A��\���R�Ћp8�Q�R��\���P��l���Q�ҡp8�P�B<����\����Ћp8�Q�RLj�j��M�QP��\����ҍ�\���P������k  �p8�Q�J��\���P�ыp8�B�P��l���Q�ҡp8�H�A�� ���R�Ћp8�Q�J������P�у��UR��,����tk  h\��������j  P��,���P��0���Q��n  ��������k  ��0���jR��z  ����u��0���P�{  �������Q��0���R�E�P�n  �p8�Q�J������P�ыp8�B�Pj j�������hd�Q�҃� ������P�M��m  �p8�Q�J������P�э�0���jR�?z  ����uP�E�P������Q�z  ���M��j  ��0����j  ��,����j  ������j  �������j  ������脋  �u��}�3ۋp8���   �P(���҉E�;�������M���l  �p8�H�A��d���R�Ћp8�Q�JSj���d���h��P�у�������R�M���j  ��p8�H�A��L���R�Ћp8�Q�J��L���PV�ыp8�B�P<����L����ҋp8�Q�RLj�j���d���QP��L����ҡp8�H�A��|���R�Ћp8�Q�R��|���P��L���Q�ҡp8�P�B<����|����Ћp8�Q�RLj�j��M�QP��|����ҍ�|���P������h  P�MQ��H���R�l  ��������i  �p8�H�A��|���R�Ћp8�Q�J��L���P�ыp8�B�P������Q�ҡp8�H�A��d���R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�hX�Q�҃�$�E�P��H����<k  �p8�Q�J�E�P�у�hBF ��H���SR襭  P蟮  ����tB��H����Mh  �p8�u��H�A�U�FR�u��Ћp8�Q�Bh��V�M�Ѕ�������KSh���M��H.���M�Q� �p8�B�P�M�Q�҃���H�����g  �p8�H�A�U�R�Ѓ��u�M�Q��  V�٬  ���M��g  �M覈  �M�g  _^�   [��]�0 W���Ȭ  ��u_�V���ڗ  ����u^_Ð�p8���   ���   ���Ѕ�tP���?����p8���   �B(���Ѕ�t�p8���   �B(���Ћ��^�   _����������U��V�uW����tW���p8���   ���   ���Ѕ�tP���ϡ���p8���   �B4����P�������p8���   �B(���Ћ���u�_�   ^]� U���4Vh��h�  h�8h�  ��  ������t���Ј �N����/���3��p8�H�A�U�R�Ћp8�Q�Jj j��E�hp�P�ыp8�B�P�M�Q�ҡp8�H�Aj j��U�hd�R�Ћp8�Q�J�E�P�ыp8�B�Pj j��M�hd�Q�҃�<�E�P�M��*� � V�M�QPj �U�Rh%� �b� ���M����%� �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�҃���^��]�������U���   �}\  V����   h@���t����wd  Ph<��M��id  P�E�P�_x  ��P�M�Q�rh  ��P�U�R�eh  ���M���d  �M���d  �M���d  ��t�����d  �E�j P�4t  ����tj �M�Q�N$��9 ���ؼ�����AH���M��d  �   ^��]� �������������VW���ǩ  ����u_^Ë�跔  ǆl      ǆt      ��t	PW���&���_�   ^���������������U���<SVW���p�  ����u�p8�H�A�UR�Ѓ�3�_^[��]� �p8�Q@�B,V�Ћp8�Q���ȋBTh%� �Ћp8�Q@�E��B,V�Ћp8�Q���ȋBTh>� �Ћp8�Q���E��B��W�Ћp8�Q�J�EWP�у��������p8�M����B�PTW�ҋM��E��p8�P�BTW�Ћp8�Q�M��RP�E�h�a  �E�P��P�M���  �M��0�  j �M���  �E�P�M��z�  �M̋���  ��t,�p8�Q�Blj Vh�a  �M��Ѕ�t�M�Q�E��#�  ���p8�B�M��P�ҡp8�P�M�B�Ћ�踗  ���Ѻ���K�9�  �p8�Q�Bj ����W�Ћp8�Q�J�EWP�у��U�R���"���P�r  ���M��ab  �p8���   �Bj j����j �T�  ���M��9�  �p8�Q�J�EP�у�_^�   [��]� ������U��SW�}�م���   V�p8���   ���   ���Ѕ�tP���̜�����5U ����t]�p8���   �B����=�F u+���O �p8���   �J�QP�҃���tP���z����p8���   �B(���Ћ���u��p8���   �B4����P���G����p8���   �B(���Ћ����=���^_[]� ���V���h�  ��u3�^Ë��Y�  ��t�P��������   ^�������V���h����3�  ��t���(�  ��tP��������   ^������U���|  SVW��3��u��}����  �؉�L���;�tC�����P����  ������ c  �p8���   �Wh   ���ЉE�;�u&������f`  �M�^�  �M�V`  3�_^[��]�0 P�E�  �M�Q�\�  �����R����p8�B�Ph3�W�M�]��҅��  �I �p8�P�BhS�M�Ћp8���   P�BH�Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A��p���R�Ћp8�Q�JWj���p���h��P�ыp8�B�Px��$��p���Q�M��ҋ�p8�H�A�ލ�p����R���Ѓ�;��  �������a  �p8�Q�J��P���P�ыp8�B�PWj���P���h��Q�҃���`���P�������_  �p8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�P�B<���M��Ћp8�Q�RLj�j���P���QP�M��ҡp8�H�A�U�R�Ћp8�Q�R�E�P�M�Q�ҡp8�P�B<���M��Ћp8�Q�RLj�j��M�QP�M��ҍE�P��(�����]  �p8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�A��`���R�Ћp8�Q�J��P���P�э�(���R�EP��0���Q�Ca  ��h���M��]  P��0���R��t���P�a  ���M��]  h\��M���\  P��0���Q������R��`  ���M��]  ��0���jP��l  ����u��0���Q�m  ����t���jR�l  ����u��t���P�cm  ����t��t���jQ�l  ������  ��`����}  �� ���WR�I�  ����  P��`����~  �� �����}  �p8�P�BhW��`���3��Ѕ��_  �p8�Q�BhS��`����Ћp8���   ���BV�Ѓ�=�   �
  �p8���   �BLV�Ѓ�P�������5\  ������WQ��k  ��;���  ������R葡  ���z�  h���M��}[  P������P�M�Q�_  ���M��!\  ������R�E�P��D���Q�j_  ��D���WR�]k  ����u?P������P�������]  P��t���Q�U�R�1_  ��P��D���P�k  ���M��   3��d$ ������VQ�3�  ������R������P�M�Q��^  ��P��D����^  �M��u[  ��D���WR��j  ����t������F�T[  ��
|��Vj�����P��������\  P��t���Q�U�R�^  ��P��D���P��j  ���M��[  ������[  ��������Z  ��D�����Z  �M���Z  �������@j�M�Q�������\  P��t���R�E�P�^  ��P������Q�jj  ���M��Z  �M��Z  �������Z  �p8�B�PhCS��`����҅��������`����c{  �]��������UZ  ��t����JZ  ��0����?Z  ��(����4Z  �p8�H�A�U�CR�]��Ћp8�Q�Bh��S�M�Ѕ�������u����h����3�  ;�t���(�  ;�tP��������p8�Q�Bh3�W�M�]��Ѕ���
  �p8�Q�BhS�M�Ћp8���   P�BH�Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A������R�Ћp8�Q�JWj�������h��P�ыp8�B�Px��$������Q�M��ҋ�p8�H�A�ލ������R���Ѓ�;��E	  �p8�Q�B����V�Ћp8�Q�J�E�VP�ы]������;����{X�v  ���  ����  �p8�J@�Q,P�ҋ�p8�P���   ��Wh�  ���Ћp8�E�ǅ����   �������Q���   ������Ph�  ���ҡp8���   �������R���E���������U��\$�C\�$�C� �p8��P�����X������   �J,P��P���P�ыp8�B���   ����P���Qh�  ���ҡp8���   ���P���R���E���\$��d����C`�$�˗ �p8��p�����x������   �J,P��p���P�ыp8�B���   ����p���Qh�  ���ҡp8���   ���p���R�Ѓ�膜  ��菈  ��訅  ��;��8  ���$    ��I �p8���   �B����=�� ��  �M��w  �p8�Q@�J$�E�PS�ыp8�B���   ��Wh�  �M��ҋ�p8�P���   Wh�  �M���j ��0�������U  ��uV;��9  �������U  �p8�Q���   Ph�  �E�P�M���P�M��!V  �M��YV  �E�P��0����zY  ��   ����   ������Q�p�  ���Y�  hh��M��\U  P������R�E�P�kY  ���M�� V  ������X  �p8�Q�J������P�ыp8�B�Pj j�������hd�Q�҃�������P������]X  �p8�Q�J������P�э����R�E�P�M�Q��X  ��P��0����X  �M��mU  �M��eU  �������ZU  j �M��T  �M��U�R��0����=Y  ��t��0���j P�d  ���E���t�E� �E�t�e���M��	U  �}� ��  ������W  �p8�Q�J������P�ыp8�B�Pj j�������h��Q�҃���P���P������lU  �p8�Q�J��������P�ыp8�B�P������QV�ҡp8�P�B<���������Ћp8�Q�RLj�j�������QP�������ҡp8�H�A������R�Ћp8�Q�R������P������Q�ҡp8�P�B<���������Ћp8�Q�RLj�j��M�QP�������ҍ�����P�M��WS  �p8�Q�J������P�ыp8�B�P������Q�ҡp8�H�A��P���R�Ћp8�Q�J������P�эU�R�EP�M�Q��V  ��h\��������R  P�U�R�����P�V  ���������AS  �����jQ�b  ����u�����R�@c  ���E�P�����Q������R�fV  �p8�H�A������R�Ћp8�Q�Jj j�������hd�P�у� ������R�������oU  �p8�H�A������R�Ѝ����jQ��a  ����uGP������R��0���P�Ab  �p8�Q�B0��j h�  �M��Ћp8�Q@�J(j�E�PS�у��������CR  ������8R  �M��0R  �M��(R  ��0����R  �M��s  3��p8���   �P(���ҋ�;������������{T  �p8�H�A������R�Ћp8�Q�JWj�������h��P�у�������R������eR  ��p8�H�A�U�R�Ћp8�Q�J�E�PV�ыp8�B�P<���M��ҋp8�Q�RLj�j�������QP�M��ҡp8�H�A������R�Ћp8�Q�R������P�M�Q�ҡp8�P�B<���������Ћp8�Q�RLj�j��M�QP�������ҍ�����P�������\P  �p8�Q�J������P�ыp8�B�P�M�Q�ҡp8�H�A������R�Ћp8�Q�J������P�у�������R��P�MQ������R��S  ��P��(���P�S  ���������QP  �p8�Q�J��`���P�ыp8�B�PWj���`���hX�Q�҃���`���P��(����R  �p8�Q�J��`���P�у�hBF ��(���WR� �  P��  ����tM��(�����O  �������O  �]��p8�H�A�U�CR�]��Ћp8�Q�Bh��S�M�Ѕ�������_Wh����`��������`���Q�) �p8�B�P��`���Q�҃���(����FO  �������;O  �p8�H�A�U�R�Ѓ��M�Q�~�  ��L���R�2�  ��������O  �M��o  �M��N  _^�   [��]�0 ������U���h  SVW��3��uЉ}���  �؉]�;�tC�� ���P����  �� ����3Q  �p8���   �Wh   ���ЉE�;�u&�� ����yN  �M�qo  �M�iN  3�_^[��]�0 P�X�  �M�Q�o�  �����e���h���M��xM  P�UR��l���P�Q  ���M��N  ��l���jQ�n]  ����u��l���R�^  ����t��l���jP�E]  ������  �M��qn  ��`���WQ��  ���  P�M���n  ��`����n  �p8�B�PhW�M�3��҅��h  �p8�P�BhS�M��Ћp8���   ���BV�Ѓ�=�   �  �p8���   �BLV�Ѓ�P��X�����L  ��X���WQ�\  ��;���  ��<���R�U�  ���>�  h���M��AL  P��<���P�M�Q�PP  ���M���L  ��X���R�E�P��P���Q�.P  ��P���WR�!\  ����uJP�����P��X����fN  P��l���Q�U�R��O  ��P��P���P�E\  ���M��zL  ������   3�������VQ��  ��X���R������P�M�Q�O  ��P��P����jO  �M��2L  ��P���WR�[  ����t������F�L  ��
|��Vj�����P��X����M  P��l���Q�U�R�EO  ��P��P���P�[  ���M���K  ������K  �������K  ��P����K  �M��K  ��<����Fj�����Q��X����EM  P��l���R�E�P��N  ��P��X���Q�$[  ���M��YK  ������NK  ��X����CK  �p8�B�PhCS�M��҅�������uЋ������Y�  ;�t���N{  ;�tP��������M���k  �p8�P�Bh3�W�M�]��Ѕ��|
  �p8�Q�BhS�M�Ћp8���   P�BH�Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A������R�Ћp8�Q�JWj�������h��P�ыp8�B�Px��$������Q�M��ҋ�p8�H�A�ލ������R���Ѓ�;��6	  �p8�Q�B����V�Ћp8�Q�J�E�VP�ы]Ѓ����Zw���{X�v  ��  ���${  �p8�J@�Q,P�ҋ�p8�P���   ��Wh�  ���Ћp8�E�ǅ ���   ��(����Q���   �� ���Ph�  ���ҡp8���   ��� ���R���E�����\����U��\$�C\�$�b� �p8���������������   �J,P������P�ыp8�B���   ��������Qh�  ���ҡp8���   �������R���E����\$��d����C`�$�� �p8���������������   �J,P������P�ыp8�B���   ��������Qh�  ���ҡp8���   �������R�Ѓ�襍  ���y  ����v  ��;��>  ���$    �d$ �p8���   �B����=�� ��  �M��h  �p8�Q@�J$�E�PS�ыp8�B���   ��Wh�  �M��ҋ�p8�P���   Wh�  �M���j ��������� G  ��ud;��G  ������F  �p8�Q���   Ph�  �E�P�M���P�M��AG  �M��yG  �E�P�������J  �M��bG  �������   ����   ��<���Q肌  ���k~  hh��M��nF  P��<���R�E�P�}J  ���M��G  �� ����I  �p8�Q�J�� ���P�ыp8�B�Pj j��� ���hd�Q�҃��� ���P�� ����oI  �p8�Q�J�� ���P�э� ���R�E�P�M�Q��I  ��P�������I  �M��F  �M��wF  ��<����lF  j �M��E  �M��U�R�������OJ  ��t������j P�U  ���E���t�E� �E�t�e���M��F  �}� ��  �� ����H  �p8�Q�J��@���P�ыp8�B�Pj j���@���h��Q�҃�������P�� ����~F  �p8�Q�J��������P�ыp8�B�P������QV�ҡp8�P�B<���������Ћp8�Q�RLj�j���@���QP�������ҡp8�H�A������R�Ћp8�Q�R������P������Q�ҡp8�P�B<���������Ћp8�Q�RLj�j��M�QP�������ҍ�����P�M��iD  �p8�Q�J������P�ыp8�B�P������Q�ҡp8�H�A������R�Ћp8�Q�J��@���P�у��UR������DD  h\��������C  P�����P��<���Q��G  ���������RD  ��<���jR�S  ����u��<���P�QT  ���M�Q��<���R�E�P�zG  �p8�Q�J�����P�ыp8�B�Pj j������hd�Q�҃� �����P�M��F  �p8�Q�J�����P�э�<���jR�S  ����uCP�E�P������Q�YS  �p8�B�P0��j h�  �M��ҡp8�H@�A(j�U�RS�Ѓ��M��_C  ��<����TC  ������IC  �M��AC  �������6C  �M��.d  3��p8���   �B(���Ћ�;�������� ����E  �p8�Q�J��0���P�ыp8�B�PWj���0���h��Q�҃�������P�� ����}C  �p8�Q�J��������P�ыp8�B�P������QV�ҡp8�P�B<���������Ћp8�Q�RLj�j���0���QP�������ҡp8�H�A������R�Ћp8�Q�R������P������Q�ҡp8�P�B<���������Ћp8�Q�RLj�j��M�QP�������ҍ�����P�������eA  P�MQ������R�4E  ����������A  �p8�H�A������R�Ћp8�Q�J������P�ыp8�B�P������Q�ҡp8�H�A��0���R�Ћp8�Q�J��t���P�ыp8�B�PWj���t���hX�Q�҃�$��t���P��������C  �p8�Q�J��t���P�у�hBF ������WR�C�  P�=�  ����tB��������@  �]��p8�H�A�U�CR�]��Ћp8�Q�Bh��S�M�Ѕ�������TWh����t���������t���Q�W�  �p8�B�P��t���Q�҃��������t@  �p8�H�A�U�R�Ѓ��M�Q跅  �U�R�n�  ����l����@@  �� ����5@  �M�-a  �M�%@  _^�   [��]�0 �������U���   SVW3���}��8�  �E�;���  ��t���P��菸���p8�Q�^(SP�B�Ћp8�Q�J��t���P�у��FdP�U�R���E�='  �}�苽  �FXP�M�Q���E�9'  �}��r�  �V\R�E�P���E�:'  �}�詽  �N`Q�U�R���E�<'  �}�落  �p8�P�M���   Whdiem��='  �-  WWS�M�Q���E�'  �}�褺  �p8�B�HW����W�ыp8�B�HWS�у���L���R��莽��P�8N  ����L�������>  ��t/j ����S������L���P���Y����N$P�� ��L����   h@��M���=  Ph<���h����=  P�M�Q�Q  ��P��L���R�A  ��P�E�P�A  ����L����B>  �M��:>  ��h����/>  �M��'>  �M�j Q�|M  ����t�N$j �U�R�7 �M���=  �}��''  �^	  ���   W�E�P���E�'  �E�    �0�  �p8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�P�Rx���E�P���ҋ��p8�H�A�ߍU��RG�Ѓ���t8j h���M�����M�Q��  �p8�B�P�M�Q�҃�3�_^[��]� �q�  �E��t�p8�Q@P�B,�Ѓ���h%� �M�Q�ˉ]܍~h����P���^  �M���]  h>� �U�R�ˍ~|���P����]  �M���]  h�� �E�P�ˍ�@  ���P���]  �M��]  �p8�Q���   j hM'  ���Ѕ��q  �p8��|  �Q�R0Ph#'  ���ҡp8�P���  �R0Ph!'  ���ҡp8�P���  �R0Ph '  ���ҡp8�P���  �R0Ph"'  ���ҡp8�P���  �R0Ph$'  ���ҡp8�P���  �R0Ph%'  ���ҡp8�P���  �R0PhF'  ���ҡp8�P���  �R0PhG'  ���ҡp8�P���  �R0PhH'  ���ҡp8�P���  �R0PhI'  ���ҡp8�P���  �R0PhJ'  ���ҡp8�P���  �R0PhK'  ���ҡp8�P�B0jhM'  ���Ћp8�Q�BDWh�� ���Ѓ��̍��   W�������d���   �E�    ;�uOj h���M�����M�Q�T�  �p8�؋B�P�M�Q�]��҃����p�������W� �����f�������$����h  9��  u<j h���M�� ���E�P�@�  �p8�Q�J�E�P�у�9��  u���%�����   u/j �M���Z  �p8�B�PD�M�Qh�a  ���   �ҍM��[  j hL��M��E ���E�P�̎  �p8�Q�J�E�P�у����P���9��  u;j h ��M��	 ���U�R萎  �p8�H�A�U�R�Ѓ�9��  u���='�����   u/j �M��JZ  �p8�Q�RD�E�Ph�a  ���   �ҍM��eZ  9��  u<j h���M������E�P��  �p8�Q�J�E�P�у�9��  u���Af�����   u/j �M���Y  �p8�B�PD�M�Qh�a  ���   �ҍM���Y  j h���M������E�P衍  �p8�Q�J�E�P�у�����&���p8�B�P���   ���ҡp8�P��h  �R$P���ҡp8�P���   P�B8h N  ���Ћp8�Q�RD���   Ph�a  ���ҡp8�P�RD���   Ph�a  ���ҡp8�P�RD��  Ph�a  ���ҡp8�P�RD��  Ph�a  ���ҡp8�P�RD��,  Ph�a  ���ҋp8�Q���   P�BDh"N  ���Ћp8�Q�B���   ���Ћp8�Q��h  �R$P���ҡp8�P���   P�B8h N  ���Ћp8�Q���   P�BDh"N  ���Ѓ}�u�����   ��P�_����������p8�Q��h  �RDWP�Nh�ҡp8�P��h  �RDS�^|P���ҡp8�P�}܍FhP�BDh%� ���Ћp8�Q�BDSh>� ���ЋM��k  �p8�Q�BTh>� ��3��Ћp8�Q���B`S���Ѓ��to�p8�Q�B`S���Ћp8�Q�E�P�BT���ЋM�;�h  u�p8�Rj���t�p8�Qj �ȋB0h�a  �Ћp8�Q�B`CS���Ѓ��u��   9~d�k  j h���M��a����M�Q��  �p8�B�P�M�Q�҃���:  �E���u�M��  3�_^[��]� �M�E�P�m  j �M��5  �M�Q�M�}��9  ��u*P��L�����4  ��L���R�M��E�   �y9  ��u2����E�t�e����L����z5  �E�t�e���M��h5  ��t/j h`��M������E�P��  �p8�Q�J�E�P�у��`W��L���R���f���P�D  ������L������5  ��t"��L���P���;���P�E  ����L�����4  ��T����������j���M���4  �M��  �P�  ���ٌ���p8���   �M�Bj j��j 誉  �}���Z��'  uR�p8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�P�Rx���E�P���E�   ���E��u�E �]���t�p8�H�A�UЃ��R�]��Ѓ��} ��   j �M��T  �M�Q���   ��T  �M���T  j �M��T  �U�R���   ��T  �M���T  j �M��|T  �E�P��  �T  �M��T  j �M��[T  �M�Q��  �T  �M��T  j �M��:T  �U�R��,  �{T  �M��cT  3�P�M쉆h  ��l  ��p  ��t  � T  �E�P���   �AT  �M��)T  ���F(��P�+������`���M��h  ��'  uR�p8�Q�J�E�P�ыp8�B�Pj j��M�h��Q�ҡp8�P�Rx���EЃ�P�N(�]����E��u�E ��t�p8�H�A�UЃ��R�]��Ѓ��} ti�p8�Q�J�E�P�ыp8�B�Pj j��M�h�Q�ҍE�P���  �p8�Q�J�E�E�P�у��}u���F(��P�7������������'  uR�p8�B�P�M�Q�ҡp8�H�Aj j��U�h��R�Ћp8�Q�Rx���EЃ�P�N(�]����E��u�E ��t�p8�H�A�UЃ��R�]��Ѓ��} �L  �p8�Q@�E��J,P�у���h>� �U�R�ω}��^|�<���P���tR  �M��\R  h%� �E�P�ύ^h����P���QR  �M��9R  ���   S�M�Q���E�'  �E�    �y�  �p8�B�P�M�Q�ҡp8�H�Aj j��U�h��R�Ћp8�Q�Rx���E�P���ҋ��p8�H�A�ߍU��RG�Ѓ����E������F(��P�������\�����p8�P�BTW�Nh�Ћp8�Q�E�BTW�N|�Ћp8�Q�M�E܋BTh�a  �Ћ}���t$�p8�Qj W�ȋBlh�a  �Ѕ�tS���b����p8�Q�M܋B8Sh N  �Ћp8�Q�M�B8Sh N  �Ћp8�Q�M��F|P�BDh>� �Ћp8�Q�M��FhP�BDh%� �Ћ���d  ����������S������M�Q���\���P���F(��P������L���R���?���P�i?  ����L����{/  �M��s/  �p8���   �Bj j����j �f�  �}�]�����)'  �B  �M�Q����H��j ��p�����O  ��p���R�M�� �wP  ��u P�M���O  �E�P�M��@�[P  �E ��t�E��@t�M�����O  �� t��p�����O  �} j �M���  h��������M�Q�m�  �p8�B�P�M�Q�҃��M��-  j hp��M�������p8�H�A�U�R�Ѓ��M�Q�U�Rjj �M��.  ���p8�H�A�U�R�Ћp8�Q�J�E�P�у�����   �UR�E�P���E�*'  �E�    �K�  �}+'  u#���U���R�-  ���E��P��N  �������},'  u#���U���R�-  ���E��P�N  �������}-'  u#���U���R�\-  ���E��P�nN  �������}.'  u#���U���R�0-  ���E��P�BN  ���{����M��S-  �M��KN  �   _^[��]� hD��s����M�Q���  �p8�B�P�M�Q�҃��M��N  �   _^[��]� ��3'  ��   �M��M  �p8�H�A��t���R�Ѓ�������  �M����`M  3���~a�M�Q�URW����  �p8�E�   �E�   �P���   �E�Ph0'  �M��ҡp8���   ��U�R�Ѓ��M�QW����  G;�|�����  �M��JM  �p8�B�P��t���Q�҃��M��*M  �   _^[��]� ��4'  ��   �M��L  �p8�H�A��t���R�Ѓ�������  �M����}L  3����z����I �M�Q�URW��� �  �p8�E�   �E�    �P���   �E�Ph0'  �M��ҡp8���   ��U�R�Ѓ��M�QW���4�  G;�|�������E'  ��   �M���K  �����l�  ��3�����   �E�P�MQW���p�  �p8�B�Pth0'  �M��ҋp8���   P�B8�Ћp8����u*�E�   �E�   �Q���   �E�Ph0'  �M��ҍU��(�E�   �E�    �Q���   �E�Ph0'  �M��ҍU��p8���   �R�Ѓ��M�QW���J�  G;��A������
�  �C�����5'  ��  �M��K  �M���J  �^�ˉ]�l�  3��E����   �U�R�E�PW���o�  �p8�Q�Bth0'  �M��Ћp8���   P�B8�Ѓ����~   �p8�Q�Bth/'  �M��Ћp8���   P�BH�Ћp8�Q�J�؍E�P�ыp8�B�P�M�QS�ҡp8�P�R8���E�PW�M��ҡp8�H�A�U�R�Ћ]��G;}�4����p8�Q�B`3�S�M��Ћ������   �d$ �p8�Q�J�E�P�у��U�RW��t���P�M������p8�Q�J�E�P�ыp8�B�H����W�ыp8�B�P��t���WQ�҃��������p8�H�A��t���RC�Ћp8�Q�B`��S�M��Ћ�����\����M��]  ��轀���M�%�  �M��I  �M��I  �   _^[��]� ��6'  ��  �p8�Q@�E��J,P�у�h%� �U�R�ȉE�~h����P���HI  �M��0I  �p8�P�B`j ���E    �Ћ؃����   �p8�Q�J��t���P�ыp8�B�PP��S�M�Q����P�M��H  �M���H  ���č�t���Qh N  P�M��������n����M��H  �p8�B�P��t���Q�ҋE�p8�Q@���EP�B`���Ћ؃���^����p8�Q�BDW�}h%� ���Ћp8�Q�RD�F|Ph>� ���ҡp8�P�BXh%� ���Ћp8�Q�BXh>� ���ЋM��\  ���!���N艒  j��L���Q���)���P�C6  ������L�������&  ����  ��L���R�������j h@��M������j h ���t���������E�P�M�Q��L����E'  P��t���R�E�P��  ��P�M�Q�  P���  �p8���B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�P��t���Q�ҡp8�H�A�U�R�Ѓ�$��u��L���VQ�5  ����L�����%  �   _^[��]� ��7'  u���B���   _^[��]� ��>'  u���a���   _^[��]� ��?'  u���
j���   _^[��]� ��@'  u"���}n��j �M��#F  �U�R�Nh�gF  � �����A'  u����u���   _^[��]� ��B'  u���&{���   _^[��]� ��L'  ��  �p8�P��x  �R0P��T  hM'  ���ҡp8�P��|  �R0Ph#'  ���ҡp8�P���  �R0Ph!'  ���ҡp8�P���  �R0Ph '  ���ҡp8�P���  �R0Ph"'  ���ҡp8�P���  �R0Ph$'  ���ҡp8�P���  �R0Ph%'  ���ҡp8�P���  �R0PhF'  ���ҡp8�P���  �R0PhG'  ���ҡp8�P���  �R0PhH'  ���ҡp8�P���  �R0PhI'  ���ҡp8�P���  �R0PhJ'  ���ҡp8�P���  �R0PhK'  ����j Wh�� �*z  ���   _^[��]� ��#'  ��   3���|  ����|  �h  �������p8�Q@P�B,�Ѓ�h�� �M��Q�ύ�@  ����P���<D  �M��$D  �p8��|  �B�P0Qh#'  ��T  �ҡp8�P�BDSh�� ���Ћ�|  Qjh#'  ���
�  �   _^[��]� ��!'  ��   3҃��  ���  ��g  ���`����p8�Q@P�B,�Ѓ�h�� �M��Q�ˍ�@  �G���P���C  �M��gC  �p8���  �B�P0Qh!'  ���ҡp8�P���  �R0Ph!'  ��T  �ҡp8�P�BDWh�� ���Ћ��  Qjh!'  ���2�  �   _^[��]� �� '  ��   3҃��  ���  �g  ����������������h�� �E�P�ˍ�@  �z���P���B  �M��B  �p8���  �Q�R0Ph '  ���ҡp8�P���  �R0Ph '  ��T  �ҡp8�P�BDWh�� ���Ћ��  Qjh '  ���e�  �   _^[��]� ��"'  ��   3҃��  ���  �Df  ���������������h�� �E�P�ˍ�@  ����P����A  �M���A  �p8���  �Q�R0Ph"'  ���ҡp8�P���  �R0Ph"'  ��T  �ҡp8�P�BDWh�� ���Ћ��  Qjh"'  ��蘻  �   _^[��]� ��$'  ��   3҃��  ���  �we  ����������8�����h�� �E�P�ˍ�@  �����P���A  �M�� A  �p8���  �Q�R0Ph$'  ���ҡp8�P���  �R0Ph$'  ��T  �ҡp8�P�BDWh�� ���Ћ��  Qjh$'  ���˺  �   _^[��]� ��%'  ��   3҃��  ���  �d  ���!������k�����h�� �E�P�ˍ�@  ����P���K@  �M��3@  �p8���  �Q�R0Ph%'  ���ҡp8�P���  �R0Ph%'  ��T  �ҡp8�P�BDWh�� ���Ћ��  Qjh%'  �����  �   _^[��]� ��F'  ��   3҃��  ���  ��c  ���T�����������h�� �E�P�ˍ�@  �F���P���~?  �M��f?  �p8���  �Q�R0PhF'  ���ҡp8�P���  �R0PhF'  ��T  �ҡp8�P�BDWh�� ���Ћ��  QjhF'  ���1�  �   _^[��]� ��G'  ��   3҃��  ���  �c  ����������������h�� �E�P�ˍ�@  �y���P���>  �M��>  �p8���  �Q�R0PhG'  ���ҡp8�P���  �R0PhG'  ��T  �ҡp8�P�BDWh�� ���Ћ��  QjhG'  ���d�  �   _^[��]� ��H'  ��   3҃��  ���  �Cb  ���������������h�� �E�P�ˍ�@  ����P����=  �M���=  �p8���  �Q�R0PhH'  ���ҡp8�P���  �R0PhH'  ��T  �ҡp8�P�BDWh�� ���Ћ��  QjhH'  ��藷  �   _^[��]� ��I'  ��   3҃��  ���  �va  ����������7�����h�� �E�P�ˍ�@  �����P���=  �M���<  �p8���  �Q�R0PhI'  ���ҡp8�P���  �R0PhI'  ��T  �ҡp8�P�BDWh�� ���Ћ��  QjhI'  ���ʶ  �   _^[��]� ��J'  ��   3҃��  ���  �`  ��� ������j�����h�� �E�P�ˍ�@  ����P���J<  �M��2<  �p8���  �Q�R0PhJ'  ���ҡp8�P���  �R0PhJ'  ��T  �ҡp8�P�BDWh�� ���Ћ��  QjhJ'  �����  �   _^[��]� ��K'  ��   3҃��  ���  ��_  ���S�����������h�� �E�P�ˍ�@  �E���P���};  �M��e;  �p8���  �Q�R0PhK'  ���ҡp8�P���  �R0PhK'  ��T  �ҡp8�P�BDWh�� ���Ћ��  QjhK'  ���0�  �   _^[��]� ��C'  ��   ��L���R�-  ��h��M��
  Ph��M���  P��L���P�M�Q�  ��P�U�R��  ���M��  �M��  �M��  j h���t���������t���P�M��  �p8�Q�J��t���P�эU�j R�(  ����u�E�P�*  ���M��&  ��L����  �   _^[��]� ��D'  ��   j h���M��2���j h����t���� ����F�M�Qj0j j�j����U��$R����P��t���P�M�Q�  ��(P�U�R��   P�^�  �p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�A��t���R�Ћp8�Q�J�E�P�у�$_^�   [��]� ��V��V�  ���    ^�������������U��V��������Et	V��A  ����^]� ���������������U��V��N�������;: �Et	V�A  ����^]� �����U��p8�H�QV�uV�ҡp8�H�U�AVR�Ћp8�Q�B<�����Ћp8�Q�M�RLj�j�QP���ҋ�^]���������U��V�u���R  �EP���W  �p8�Q�J�EP�у���^]� �����������U���X�E$jP�_&  ����uS�p8�Q�J�E�VP�ыp8�B�Pj j��M�hP�Q�ҍE�P�@�  �p8�Q�J���E�P�у���^tY�U$R�&  ����ua�p8�H�A�U�R�Ћp8�Q�Jj j��E�h �P�эU�R��  �p8�H�A�U�R�Ѓ��M�C  �M$�;  3���]�8 �#  j �MQ�ȉE���#  �M���tq�$  ��th�M��U�R�$  �E�P�MQ�U�R�Q  �E�P�M$Q�U�R�@  j�E�P�M�Q�%  ��$�Mą�tO��  �M��  �M��  �M��#  ��u��E�P�m#  ���M�E�    �  �M$�  �   ��]�8 �s  �M��k  �M��c  �U�R�*#  ���E�    � ��������������U���0  �}vF VW���M  �u���B  �>�  �6  �JZ  ���)  ��P���P�6Z  ���L  �M�Q�&Z  ���OK  �U�R��P���P������Q�(  ���M��M  �U�R�M���  j h���M�������E�P�M�Q�U�R������p8�H�A�U�R�ЍU���R���������P�����������Q��P���R��l���P�  ����V�M���  V��������  �M��  j h���M��[����M�Q��@���R�M���  P�E�P�N����p8�Q�J��@���P�ыp8�B�P�M�Q�҃��E���P�������$���Q���k���������R�������  ��t?��l���jP��"  ����u)����$�����R�>  ����l�����P�-  ���V�����$����[  �p8�Q�J�E�P�у��������;  �M��3  ��l����(  ������  �p8�B�P�M�Q�ҡp8�H�A�U�R�Ѓ���������  �M���  ��P�����  _�   ^��]� ������������U��p8�H�A���U�VR�Ћp8�Q�Jj j��E�h��P��j j h�  h@8h    �U�Rhϗ �X ��p8�H�A�U�R�Ѓ�4��^��]����������������U��V���4 �Et	V��;  ����^]� ���������������Vh0�jh�8j�<  ������t���L4 �����^�3�^���������������U��E��u�`8�MP�EPQ��  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h��j;h�8j��;  ����t
W���  �3��F��u_^]� �~ t3�9_��^]� �p8�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   �p8�H<�Q��3Ʌ����^��������������̃y t�   ËA��uËp8�R<P��JP�у��������U����u�p8�H�]� �p8�J<�URP�A�Ѓ�]� ���������������U��`8��u�p8�H�]Ëp8�J<�URP�A�Ѓ�]�U��`8��$V��u�p8�H�1��p8�J<�URP�A�Ѓ����p8�Q�J�E�SP�ыp8�B�P�M�QV�ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@�� j �M�Q�U�R�M��Ћp8�Q�J���E�P���у���[t.�p8�B�u�HV�ыp8�B�P�M�Q�҃���^��]áp8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�u�QV�ҡp8�H�A�U�VR�Ћp8�Q�J�E�P�у���^��]���������������U��`8��$SV��u�p8�H�1��p8�J<�URP�A�Ѓ����p8�Q�J�E�P�ыp8�B�P�M�QV�ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@�� j �M�Q�U�R�M��Ћp8�Q�J���E�P���у���t/�p8�B�u�HV�ыp8�B�P�M�Q�҃���^[��]áp8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@��j �M�Q�U�R�M��Ћp8�Q�J���E�P���у����3����p8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�u�QV�ҡp8�H�A�U�VR�Ћp8�Q�J�E�P�у���^[��]����������������U��`8��$SV��u�p8�H�1��p8�J<�URP�A�Ѓ����p8�Q�J�E�P�ыp8�B�P�M�QV�ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@�� j �M�Q�U�R�M��Ћp8�Q�J���E�P���у���t/�p8�B�u�HV�ыp8�B�P�M�Q�҃���^[��]áp8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@��j �M�Q�U�R�M��Ћp8�Q�J���E�P���у����3����p8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@��j �M�Q�U�R�M��Ћp8�Q�J���E�P���у���������p8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҋu�E�P���c����p8�Q�J�E�P�у���^[��]�������U��`8��$SV��u�p8�H�1��p8�J<�URP�A�Ѓ����p8�Q�J�E�P�ыp8�B�P�M�QV�ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@�� j �M�Q�U�R�M��Ћp8�Q�J���E�P���у���t/�p8�B�u�HV�ыp8�B�P�M�Q�҃���^[��]áp8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@��j �M�Q�U�R�M��Ћp8�Q�J���E�P���у����3����p8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M��ҡp8�H�A�U�R�Ћp8�Q�Jj j��E�h��P�ыp8�B�@@��j �M�Q�U�R�M��Ћp8�Q�J���E�P���у���������p8�P�E��RHjP�M��ҡp8�P�E�M��RLj�j�PQ�M���j h���M������p8�P�R@j �E�P�M�Q�M��҅��p8�H�A�U�R���Ѓ���t/�p8�Q�u�BV�Ћp8�Q�J�E�P�у���^[��]Ëp8�M��B�PHjQ�M��ҡp8�P�E�M��RLj�j�PQ�M��ҋu�E�P���+����p8�Q�J�E�P�у���^[��]���������������U��p8�H<�A]����������������̡p8�H<�Q�����V��~ u>���t�p8�Q<P�B�Ѓ��    W�~��t���  W�T0  ���F    _^��������U���V�E�P���  ��P��������M���I  ��^��]��̃=h8 uK�`8��t�p8�Q<P�B�Ѓ��`8    �l8��tV���   V��/  ���l8    ^������������U���8�p8�H�AS�U�V3�R�]��Ћp8�Q�JSj��E�h��P�ыp8�B<�P�M�Q�ҋ�p8�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��M �M�Q�U�R�M��XM ����   W�}�}���   �p8���   �U��ATR�Ћ�����tB�p8�Q�J�E�P���у��U�Rj�E�P���\����p8�Q�ȋBxW���E���t�E� ��t�p8�Q�J�E�P����у���t�p8�B�P�M�Q����҃��}� u"�E�P�M�Q�M��L ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_�p8�H�A�U�R�Ћp8�Q�JSj��E�h��P�ыp8�B<�P�M�Q�ҋ�p8�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��K �M�Q�U�R�M���K ���p  W�}��I �E����   �p8���   �U��ATR�Ћ�������   �p8�Q�J�E�P���ыp8�B���   ���M�Qj�U�R���Ћp8�Q�J���E�P�ыp8�B�P�M�QV�ҡp8�H�A�U�R�Ћp8�Q�Bx��W�M����E��t�E ��t�p8�Q�J�E�P����у���t�p8�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�p8���   P�BH�Ћp8�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��rJ ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M���I �EP�M�Q�M�u��u�J ����   �u���E���tA��t<��uZ�p8���   �M�PHQ�ҋp8�Q���ȋBxV�Ѕ�u-�   ^��]Ëp8���   �E�JTP��VP�[�������uӍUR�E�P�M��I ��u�3�^��]����������V��~ u>���t�p8�Q<P�B�Ѓ��    W�~��t���J  W�+  ���F    _^��������U��E�p8� ]��U��p8�P�EP�EP�EPQ�J�у�]� �����������̡p8V��H�QV�ҡp8�H$�QDV�҃���^�����������U��p8V��H�QV�ҡp8�H$�QDV�ҡp8�U�H$�AdRV�Ѓ���^]� ��U��p8V��H�QV�ҡp8�H$�QDV�ҡp8�U�H$�ARV�Ѓ���^]� ��U��p8V��H�QV�ҡp8�H$�QDV�ҡp8�H$�U�ALVR�Ѓ���^]� �̡p8V��H$�QHV�ҡp8�H�QV�҃�^�������������U��p8�P$�EPQ�JL�у�]� ����U��p8�P$�R]�����������������U��p8�P$�Rl]����������������̡p8�P$�Bp����̡p8�P$�BQ�Ѓ����������������U��p8�P$��VWQ�J�E�P�ыp8�u���B�HV�ыp8�B�HVW�ыp8�B�P�M�Q�҃�_��^��]� ���U��p8�P$�EPQ�J�у�]� ����U��p8�P$��VWQ�J �E�P�ыp8�u���B�HV�ыp8�B$�HDV�ыp8�B$�HLVW�ыp8�B$�PH�M�Q�ҡp8�H�A�U�R�Ѓ� _��^��]� ���U��p8�P$��VWQ�J$�E�P�ыp8�u���B�HV�ыp8�B$�HDV�ыp8�B$�HLVW�ыp8�B$�PH�M�Q�ҡp8�H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e����p8�Q$�JH�E�P�ыp8�B�P�M�Q�҃���^��]� ����̡p8�P$�B(Q��Yáp8�P$�BhQ��Y�U��p8�P$�EPQ�J,�у�]� ����U��p8�P$�EPQ�J0�у�]� ����U��p8�P$�EPQ�J4�у�]� ����U��p8�P$�EPQ�J8�у�]� ����U��p8�UV��H$�ALVR�Ѓ���^]� ��������������U��p8�H�QV�uV�ҡp8�H$�QDV�ҡp8�H$�U�ALVR�Ћp8�E�Q$�J@PV�у���^]�U��p8�UV��H$�A@RV�Ѓ���^]� ��������������U��p8�P$�EPQ�J<�у�]� ����U��p8�P$�EPQ�J<�у����@]� ���������������U��p8�P$�EP�EPQ�JP�у�]� U��p8�P$�EPQ�JT�у�]� ���̡p8�H$�QX�����U��p8�H$�A\]�����������������U��p8�P$�EP�EP�EPQ�J`�у�]� �����������̡p8�H(�������U��p8�H(�AV�u�R�Ѓ��    ^]��������������U��p8�P(�R]����������������̡p8�P(�B�����U��p8�P(�R]�����������������U��p8�P(�R]�����������������U��p8�P(�R ]�����������������U��p8�P(�E�RjP�EP��]� ��U��p8�P(�E�R$P�EP�EP��]� �p8�P(�B(����̡p8�P(�B,����̡p8�P(�B0�����U��p8�P(�R4]�����������������U��p8�P(�RX]�����������������U��p8�P(�R\]�����������������U��p8�P(�R`]�����������������U��p8�P(�Rd]�����������������U��p8�P(�Rh]�����������������U��p8�P(�Rx]�����������������U��p8�P(�Rl]�����������������U��p8�P(�Rt]�����������������U��p8�P(�Rp]�����������������U��p8�P(�BpVW�}W���Ѕ�t:�p8�Q(�Rp�GP���҅�t"�p8�P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U��p8�P(�BtVW�}W���Ѕ�t:�p8�Q(�Rt�GP���҅�t"�p8�P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U����p8�E�    �E�    �P(�RhV�E�P���҅���   �E���uG�p8�H�A�U�R�Ћp8�Q�E�RP�M�Q�ҡp8�H�A�U�R�Ѓ��   ^��]� �p8�Qh��h`  P���   �Ћp8���E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P��  ��3�^��]� �M��U�j IQ�MR�����E�P�  ���   ^��]� ���������������U��p8��V��H�A�U�R�Ѓ��M�Q������^��u�p8�B�P�M�Q�҃�3���]� �p8�H$�E�I�U�RP�ыp8�B�P�M�Q�҃��   ��]� �U��Q�p8�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U��p8�P(�R8]�����������������U��p8�P(�R<]�����������������U��p8�P(�R@]�����������������U��p8�P(�RD]�����������������U��p8�P(�RH]�����������������U��p8�P(�E�R|P�EP��]� ����U��p8�P(�RL]�����������������U��p8�E�P(�BT���$��]� ���U��p8�E�P(�BPQ�$��]� ����̡p8�H(�Q�����U��p8�H(�AV�u�R�Ѓ��    ^]��������������U��p8�P(���   ]��������������U��p8�H(�A]����������������̡p8�H,�Q,����̡p8�P,�B4�����U��p8�H,�A0V�u�R�Ѓ��    ^]�������������̡p8�P,�B8�����U��p8�P,�R<��VW�E�P�ҋu���p8�H�QV�ҡp8�H$�QDV�ҡp8�H$�QLVW�ҡp8�H$�AH�U�R�Ћp8�Q�J�E�P�у�_��^��]� �������U��p8�P,�E�R@��VWP�E�P�ҋu���p8�H�QV�ҡp8�H�QVW�ҡp8�H�A�U�R�Ѓ�_��^��]� ��̡p8�H,�j j �҃��������������U��p8�P,�EP�EPQ�J�у�]� U��p8�H,�AV�u�R�Ѓ��    ^]�������������̡p8�P,�B����̡p8�P,�B����̡p8�P,�B����̡p8�P,�B ����̡p8�P,�B$����̡p8�P,�B(�����U��p8�P,�R]�����������������U��p8�P,�R��VW�E�P�ҋu���p8�H�QV�ҡp8�H$�QDV�ҡp8�H$�QLVW�ҡp8�H$�AH�U�R�Ћp8�Q�J�E�P�у�_��^��]� �������U��p8�H��D  ]��������������U��p8�H��H  ]��������������U��p8�H��L  ]��������������U��p8�H�I]�����������������U��p8�H�A]�����������������U��p8�H�I]�����������������U��p8�H�A]�����������������U��p8�H�I]�����������������U��p8�H���  ]��������������U��p8�H�A]�����������������U���V�u�E�P��������p8�Q$�J�E�P�у���u-�p8�B$�PH�M�Q�ҡp8�H�A�U�R�Ѓ�3�^��]Ëp8�Q�J�E�jP�у���u=�U�R��������u-�p8�H$�AH�U�R�Ћp8�Q�J�E�P�у�3�^��]Ëp8�B�HjV�у���u�p8�B�HV�у����I����p8�Q$�JH�E�P�ыp8�B�P�M�Q�҃��   ^��]�����������U��p8�H�A ]�����������������U��p8�H�I(]�����������������U��p8�H��  ]��������������U��p8�H��   ]��������������U��p8�H��  ]��������������U��p8�H��  ]��������������U��p8�H�A$��V�U�WR�Ћp8�Q�u���BV�Ћp8�Q$�BDV�Ћp8�Q$�BLVW�Ћp8�Q$�JH�E�P�ыp8�B�P�M�Q�҃�_��^��]������U��p8�H���  ��V�U�WR�Ћp8�Q�u���BV�Ћp8�Q$�BDV�Ћp8�Q$�BLVW�Ћp8�Q$�JH�E�P�ыp8�B�P�M�Q�҃�_��^��]���U��p8�H���  ]��������������U���<��8SVW�E�    ��t�E�P�   ��������/�p8�Q�J�E�P�   �ыp8�B$�PD�M�Q�҃��}�p8�H�u�QV�ҡp8�H$�QDV�ҡp8�H$�QLVW�҃���t)�p8�H$�AH�U�R����Ћp8�Q�J�E�P�у���t&�p8�B$�PH�M�Q�ҡp8�H�A�U�R�Ѓ�_��^[��]���U��p8�H�U���  ��VWR�E�P�ыp8�u���B�HV�ыp8�B$�HDV�ыp8�B$�HLVW�ыp8�B$�PH�M�Q�ҡp8�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡p8�H���   ��U��p8�H���   V�uV�҃��    ^]�������������U��p8�P�]��p8�P�B����̡p8�P���   ��U��p8�P�R`]�����������������U��p8�P�Rd]�����������������U��p8�P�Rh]�����������������U��p8�P�Rl]�����������������U��p8�P�Rp]�����������������U��p8�P�Rt]�����������������U��p8�P���   ]��������������U��p8�P�Rx]�����������������U��p8�P���   ]��������������U��p8�P�R|]�����������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P�EPQ��  �у�]� �U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��E��t �p8�R P�B$Q�Ѓ���t	�   ]� 3�]� U��p8�P �E�RLQ�MPQ�҃�]� U��E��u]� �p8�R P�B(Q�Ѓ��   ]� ������U��p8�P�R]�����������������U��p8�P�R]�����������������U��p8�P�R]�����������������U��p8�P�R]�����������������U��p8�P�R]�����������������U��p8�P�R]�����������������U��p8�P�E�R\P�EP��]� ����U��p8�E�P�B ���$��]� ���U��p8�E�P�B$Q�$��]� �����U��p8�E�P�B(���$��]� ���U��p8�P�R,]�����������������U��p8�P�R0]�����������������U��p8�P�R4]�����������������U��p8�P�R8]�����������������U��p8�P�R<]�����������������U��p8�P�R@]�����������������U��p8�P�RD]�����������������U��p8�P�RH]�����������������U��p8�P�RL]�����������������U��p8�P�RP]�����������������U��p8�P���   ]��������������U��p8�P�RT]�����������������U��p8�P�EPQ��  �у�]� �U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P�RX]����������������̡p8�P���   ��U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]��������������U��p8�P���   ]�������������̡p8�P���   ��U��p8�P���   ]�������������̡p8�P���   ��p8�P���   ��p8�P���   ��U��p8�H���   ]��������������U��p8�H��   ]��������������U��p8�H�U�E��VWRP���  �U�R�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�_��^��]������������U��p8�H���  ]��������������U��p8�P(�BPVW�}�Q�]���E�$�Ѕ�tM�p8�G�Q(�]�E�BPQ���$�Ѕ�t,�p8�G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U��p8�P(�BTVW�}����$���Ѕ�tE�p8�G�Q(�BT�����$�Ѕ�t(�p8�G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U��p8�P(�} �R8����P��]� �U��p8�P�BdS�]VW��j ���Ћp8�Q�����   h��Fh�  V�Ћp8���E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћp8�Q(�BHV���Ѕ�t �p8�Q(�E�R VP���҅�t�   �3��EP�B  ��_��^[]� ������U���V�E���MP�K���P���#����p8�Q�J���E�P�у���^��]� ��̡p8�P�BVj j����Ћ�^���������U��p8�P�E�RVj P���ҋ�^]� U��p8�P�E�RVPj����ҋ�^]� �p8�P�B�����U��p8�P���   Vj ��Mj V�Ћ�^]� �����������U��p8�P�EPQ�J�у�]� ����U��p8�P�EPQ�J�у����@]� ���������������U��p8�P�E�RtP�ҋp8���   P�BX�Ѓ�]� ���U��p8�P�E�Rlh#  P�EP��]� ���������������U��p8�P�E�RlhF  P�EP��]� ���������������U��p8�P�E�RtP�ҋp8���   �M�R`QP�҃�]� ���������������U��p8�P���   ]��������������U��p8�P�E���   P�҅�u]� �p8���   P�B�Ѓ�]� ��������U��M��P]����U��M��P]����U��M��P]����V���4��F    �p8�HP�h0mVh mhm�҉F����^����������̃y �4�u�p8�PP�A�JP��Y��U��A��u]� �p8�QP�M�Rj Q�MQP�҃�]� ��U��A��t�p8�QP�M�RQP�҃�]� ������������U��A��t�p8�QP�M�RQP�҃�]� �����������̡p8�HP���   ��U��p8�HP���   ]�������������̡p8�HP�QP�����U��p8�HP�AT]����������������̋��     �@    �V����t)�p8�QPP�BL�Ћp8�QP��J<P�у��    ^�������������U��SV�ً3�W;�t�p8�QPP�B<�Ѓ��3�s�}�Eh0mW�C�p8�QP�J8h mhmP�EP�у�9u�~M�I ���z u!���@   �p8�QP���H�RQ�҃��p8�HP��A@VR�Ћ�F��;u�A|�3�9_^��[]� ��������U��SVW��3�9w~<�]�p8�HP��A@VR�Ѓ���t-�p8�QPj SjP�B�Ѓ���tF;w|�_^�   []� �p8�QP��JLP�у�_^3�[]� �����������̡p8�PP��JDP�у�������������̡p8�PP��JHP��Y��������������̡p8�PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ �4�u�p8�HP�V�AR�Ѓ��Et	V�N  ����^]� ����U��V�u���t�p8�QP��Ѓ��    ^]���������̡p8�H��@  hﾭ���Y����������U��E��t�p8�QP��@  �Ѓ�]����������������U��p8�H���  ]��������������U��p8�H��  ]�������������̡p8�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�6� ������u_^]Ã} tWj V�� ��_������F�t8   ^]���U��p8�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW躆 ������u_^]�Wj V�v� ��_������F�t8   ^]�������������U��p8�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�:� ������u_^]�Wj V��� ��_������F�t8   ^]�������������U��p8�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW躅 ������u_^]�Wj V�v� ��_������F�t8   ^]�������������U��p8�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�:� ������u_^]�Wj V��� ��_������F�t8   ^]�������������U��M��t-�=t8 t�y���A�uP�(� ��]áp8�P�Q�Ѓ�]��������U��M��t-�=t8 t�y���A�uP�� ��]áp8�P�Q�Ѓ�]��������U��p8�H�U�R�Ѓ�]���������U��p8�H�U�R�Ѓ�]���������U��p8�E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��� ������u_^]�Wj V貄 ��_������F�t8   ^]���������U��p8�E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   �p8��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�� ������u_^]�Wj V�Ã ��_������F�t8   ^]����������U��E��w�   �p8��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�t� ������u_^]�Wj V�0� ��_������F�t8   ^]�������U��p8�H�U�R�Ѓ�]���������U��p8�H�U�R�Ѓ�]���������U��p8�H�U�R�Ѓ�]���������U��p8�H�U�R�Ѓ�]���������U��p8�Hp�]��p8�Hp�h   �҃�������������U��V�u���t�p8�QpP�B�Ѓ��    ^]���������U��p8�Pp�EP�EPQ�J�у�]� U��p8�Pp�EP�EPQ�J�у�]� U��p8�Pp�EP�EPQ�J�у�]� U��p8�Pp�EPQ�J�у�]� ���̡p8�HL���   ��U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�HL�������U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�PL���   Q�Ѓ�������������U��p8�PL�EP�EPQ���   �у�]� �������������U��p8V��HL���   V�҃���u�p8�U�HL���   j RV�Ѓ�^]� �p8���   �ȋBP�Ћp8���   �MP�BH��^]� �����̡p8�PL��(  Q�Ѓ�������������U��p8�PL�EP�EPQ��,  �у�]� ������������̡p8�HL�Q�����U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�PL�E�R��VPQ�M�Q�ҋu��P��������M�������^��]� ����U��p8�PL�EPQ���   �у�]� �U��p8�PL�EP�EPQ�J�у�]� �p8�PL�BQ�Ѓ���������������̡p8�PL�BQ�Ѓ���������������̡p8�PL�BQ�Ѓ����������������U��p8�PL�EP�EP�EPQ�J �у�]� ������������U��p8�PL�EPQ��4  �у�]� �U��p8�PL�EP�EP�EPQ�J$�у�]� ������������U��p8�PL�EP�EP�EP�EPQ�J(�у�]� �������̡p8�PL�B,Q�Ѓ���������������̡p8�PL�B0Q�Ѓ����������������U��p8�PL�EP�EPQ��  �у�]� ������������̡p8�PL���   Q�Ѓ�������������U��p8�PL�E��  ��VPQ�M�Q�ҋu��P��������M��������^��]� ̡p8�PL�B4Q�Ѓ���������������̡p8�PL�B8j Q�Ѓ��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL���   ]��������������U��p8�PL�EPQ�J<�у�]� ���̡p8�PL�BQ��Y�U��p8�PL�EP�EPQ�J@�у�]� U��p8�PL�Ej PQ�JD�у�]� ��U��p8�PL�Ej PQ�JH�у�]� ��U��p8�PL�EjPQ�JD�у�]� ��U��p8�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�贰  W�M�Q�U�R���t�  ���M�����  ��t�p8���   ��U�R�Ѓ�_^3�[��]Ëp8���   �J8�E�P�ыp8�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ���  j�M�Q�U�R�����  �M��e�  �p8���   ��U�R�Ѓ�^��]�����������U���$�p8�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��z�  j�E�P�M�Q���Y�  �M���  �p8���   ��M�Q�҃�_^��]� ��U���$�p8�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}����  j�E�P�M�Q�����  �M��a�  �p8���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�蔮  W�M�Q�U�R���T�  ���M������  ��t+�u���I����p8���   ��U�R�Ѓ�_��^[��]� �p8���   �JL�E�P�ыu��P�������p8���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��ԭ  W�M�Q�U�R����  ���M����7�  ��t+�u�������p8���   ��U�R�Ѓ�_��^[��]� �p8���   �JL�E�P�ыu��P��������p8���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���  W�M�Q�U�R�����  ���M����w�  _^��[t�p8���   ��U�R�������]Ëp8���   �J<�E�P���]��p8���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��d�  W�M�Q�U�R���$�  ���M����Ǟ  ��t�p8���   ��U�R�Ѓ�_^3�[��]Ëp8���   �J8�E�P�ыp8�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}�贫  W�M�Q�U�R���t�  ���M�����  ��t-��u�p8����   ���^�U�R�Ѓ�_��^[��]� �p8���   �JP�E�P�ы�u�H��P�@�N�p8�V���   �
�F�E�P�у�_��^[��]� �����̡p8�PL���   Q��Y��������������U��p8�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U��p8�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��$�  W�M�Q�U�R�����  ���M���臜  ��t-��u�p8����   ���^�U�R�Ѓ�_��^[��]� �p8���   �JP�E�P�ы�u�H��P�@�N�p8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��T�  W�M�Q�U�R����  ���M���跛  ��t-��u�p8����   ���^�U�R�Ѓ�_��^[��]� �p8���   �JP�E�P�ы�u�H��P�@�N�p8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�脨  W�M�Q�U�R���D�  ���M�����  ��t-��u�p8����   ���^�U�R�Ѓ�_��^[��]� �p8���   �JP�E�P�ы�u�H��P�@�N�p8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�货  W�M�Q�U�R���t�  ���M�����  ��t�p8���   ��U�R�Ѓ�_^3�[��]Ëp8���   �J8�E�P�ыp8�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ���  j�M�Q�UR�����  �M�f�  �p8���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�菦  j�U�R�E�P���n�  �M����  �p8���   �
�E�P�у�^��]� ��������U���$�p8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
�  j�E�P�M�Q�����  �M��q�  �p8���   ��M�Q�҃�_^��]� ��U���$�p8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}�芥  j�E�P�M�Q���i�  �M���  �p8���   ��M�Q�҃�_^��]� ��U���$�p8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
�  j�E�P�M�Q�����  �M��q�  �p8���   ��M�Q�҃�_^��]� ��U���$�p8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}�芤  j�E�P�M�Q���i�  �M���  �p8���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���  j�U�R�E�P�����  �M�膖  �p8���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}�责  W�M�Q�U�R���t�  ���M�����  ��t-��u�p8����   ���^�U�R�Ѓ�_��^[��]� �p8���   �JP�E�P�ы�u�H��P�@�N�p8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���  W�M�Q�U�R����  ���M����G�  ��t�p8���   ��U�R�Ѓ�_^3�[��]Ëp8���   �J8�E�P�ыp8�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��4�  W�M�Q�U�R�����  ���M���藔  ��t�p8���   ��U�R�Ѓ�_^3�[��]Ëp8���   �J8�E�P�ыp8�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$�p8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J�  j�E�P�M�Q���)�  �M�豓  �p8���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��ߠ  j�U�R�E�P����  �M��F�  �p8���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��o�  j�U�R�E�P���N�  �M��֒  �p8���   �
�E�P�у�^��]� ��������U��p8�H���   ]��������������U��p8�H���   ]�������������̡p8�H���   ��p8�H���   ��U��p8�H���   V�u�R�Ѓ��    ^]�����������U��p8�H���   ]��������������U��p8�HL�QV�ҋ���u^]áp8�H�U�ER�UP���  RV�Ѓ���u�p8�Q@�BV�Ѓ�3���^]����������U��p8�H�U�E���  R�U�� P�ERP�у�]������U��p8�H���   ]��������������U��p8�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡p8�PL�BLQ�Ѓ���������������̡p8�PL�BPQ�Ѓ����������������U��p8�PL�EP�EPQ�JT�у�]� U��p8�PL�EPQ��  �у�]� �U��p8�PL�EPQ���   �у�]� ̡p8�PL�BXQ�Ѓ����������������U��p8�PL�EP�EP�EPQ�J\�у�]� ������������U���4�p8SV��HL�QW�ҋ�3ۉ}�;��x  �M�������p8�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡp8���   �BSSW���Ѕ���   �p8�QL�BW�Ћ���;���   ��    �p8���   �B(���ЍM�Qh�   ���u��  ������   �M�;���   �p8���   ���   S��;�tm�p8���   �ȋB<V�Ћp8���   ���   �E�P�у�;�t�p8�B@�HV�у���;��\����}��M���   �M�������_^[��]� �}��p8�B@�HW�ыp8���   ���   �M�Q�҃��M��   �M������_^3�[��]� �����̡p8�PL�B`Q�Ѓ���������������̡p8�PL�BdQ�Ѓ����������������U��p8�PL�EPQ�Jh�у�]� ���̡p8�PL��D  Q�Ѓ������������̡p8�PL�BlQ�Ѓ����������������U��p8�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh��h��h`�hP�R�Q�U R�UR�UR�U���A�$�5p8�vLRP���   Q�Ѓ�4^]�  ������̡p8�PL���   Q�Ѓ�������������U��p8�PL�EP�EP�EPQ��   �у�]� ���������U��p8�PL��H  ]�������������̡p8�PL��L  ��U��p8�PL��P  ]��������������U��p8�PL��T  ]��������������U��p8�PL�EP�EP�EP�EP�EPQ���   �у�]� �U��p8�PL�EP�EP�EPQ���   �у�]� ���������U��p8�PL�EP�EP�EP�EPQ��   �у�]� �����U��p8�HL���   ]��������������U��p8�HL���   ]��������������U��p8�HL���   ]�������������̡p8�HL��  ��p8�HL��@  ��h�8Ph^� � �  ���������������U��Vh�8j\h^� �����  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� �p8V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�p8�QLjP���   ���ЋM��U�Rh=���M�}��  ���p8���   ���   �U�R�Ѓ��M��u��<  ��_^��]Ëp8���   ���   �E�P�у��M��u��  _�   ^��]����U��� �p8V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�p8�QLjP���   ���ЋM��U�Rh<���M�}��3  ���p8���   ���   �U�R�Ѓ��M��u��l  ��_^��]Ëp8���   ���   �E�P�у��M��u��>  _�   ^��]���̡p8V�񋈈   ���   V�҃��    ^���������������U��p8�P8�EPQ�JD�у�]� ���̡p8�H8�Q<�����U��p8�H8�A@V�u�R�Ѓ��    ^]�������������̡p8�H8�������U��p8�H8�AV�u�R�Ѓ��    ^]��������������U��p8�P8�EP�EP�EPQ�J�у�]� ������������U��p8�P8�EP�EPQ�J�у�]� �p8�P8�BQ�Ѓ����������������U��p8�P8�EPQ�J �у�]� ����U��p8�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U��p8�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U��p8�P8�EP�EPQ�J(�у�]� U��p8�P8�EP�EP�EPQ�J,�у�]� ������������U��p8�P8�EP�EP�EPQ�J�у�]� ������������U��p8�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U��p8�P8�EP�EPQ�J0�у�]� U��p8�P8�EP�EP�EPQ�J4�у�]� ������������U��p8�P8�EPQ�J8�у�]� ����U��p8�H��x  ]��������������U��p8�H��|  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H�A,]�����������������U��p8�H�QV�uV�ҡp8�H�Q8V�҃���^]�����̡p8�H�Q<�����U��p8�H�I@]����������������̡p8�H�QD����̡p8�H�QH�����U��p8�H�AL]�����������������U��p8�H�IP]�����������������U��p8�H��<  ]��������������U��p8�H��,  ]��������������U��p8�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡p8�H���   ��p8�H���  ��U��p8�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U��p8�H�A]�����������������U��p8�H��\  ]��������������U��p8�H�AT]�����������������U��p8�H�AX]�����������������U��p8�H�A\]����������������̡p8�H�Q`����̡p8�H�Qd����̡p8�H�Qh�����U��p8�H�Al]�����������������U��p8�H�Ap]�����������������U��p8�H�At]�����������������U��p8�H��D  ]��������������U��p8�H��  ]��������������U��p8�H�Ix]�����������������U��p8�H��@  ]��������������U��V�u���r����p8�H�U�A|VR�Ѓ���^]���������U��p8�H���   ]��������������U��p8�H��h  ]��������������U��p8�H��d  ]��������������U��p8�H���  ]�������������̡p8�H���   ��U��p8�H��l  ]��������������U��p8�H��   ]��������������U��p8�H��  ]��������������U��V�u��������p8�H���   V�҃���^]���������̡p8�H��`  ��U��p8�H��  ]��������������U��p8�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U��p8�H���  ]��������������U��U�E�p8�H�E���   R���\$�E�$P�у�]�U��p8�H���   ]��������������U��p8�H���   ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���   ]��������������U��p8�H���   ]��������������U��p8�H���   ]��������������U��p8�H���   ]��������������U��p8�H���   ]��������������U��p8�H���   ]��������������U��p8�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��p8�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��p8�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��p8�H��8  ]��������������U��V�u(V�u$�E�@�p8�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@�p8�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��p8�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U��p8�P0�EP�EP�EP�EPQ���   �у�]� ����̡p8�P0���   Q�Ѓ�������������U��p8�P0�EP�EPQ���   �у�]� �������������U��p8�P0�EP�EP�EP�EPQ���   �у�]� ����̡p8�P0���   Q�Ѓ������������̡p8�H0���   ��U��p8�H0���   V�u�R�Ѓ��    ^]�����������U��p8�H��H  ]��������������U��p8�H��T  ]�������������̡p8�H��p  ��p8�H���  ��U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �p8���   �Qj PV�ҡp8���   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M��Z���P�E�hicMCP�k������M������p8���   �JT�E�P�у���u(�u��������p8���   ��M�Q�҃���^��]áp8���   �AT�U�R�Ћu��P��������p8���   �
�E�P�у���^��]�������������U��p8�H��  ]��������������U��p8�H��\  ]��������������U��p8�H�U��t  ��V�uVR�E�P�у����C����M��{�����^��]�����U��p8�H�U���  ��VWR�E�P�ыp8�u���B�HV�ыp8�B�HVW�ыp8�B�P�M�Q�҃�_��^��]����������������U��p8�H�U���  ��VWR�E�P�ыp8�u���B�HV�ыp8�B�HVW�ыp8�B�P�M�Q�҃�_��^��]����������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H�U�E��VWj R�UP�ERP��t  �U�R�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�(_��^��]��U��p8�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �p8���   j P�BV�Ћp8���   �
�E�P�у�$��^��]���U��p8�H��8  ]��������������U���  �@#3ŉE��M�EPQ������h   R�1� ����|	=�  |#��p8�H��0  hD�hF  �҃��E� �p8�H��4  ������Rh���ЋM�3̓��O ��]�������U��p8�H��  ��V�U�WR�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�_��^��]����U��p8�H��  ��V�U�WR�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�_��^��]����U��p8�H��p  ��$�҅�trh���M��9����p8�P�E�R4Ph���M��ҡp8�P�E�R4Ph���M���j �E�P�M�hicMCQ�����p8���   ��M�Q�҃��M�������]�U��p8�H��p  ��$V�҅�u�p8�H�u�QV�҃���^��]�Wh!���M�茽���p8�P�E�R4Ph!���M���j �E�P�M�hicMCQ�����p8���   �QHP�ҋu���p8�H�QV�ҡp8�H�QVW�ҡp8���   ��U�R�Ѓ�$�M��M���_��^��]������U��p8�H��p  ��$V�҅�u�p8�H�u�QV�҃���^��]�Wh����M�輼���p8�P�E�R4Ph����M���j �E�P�M�hicMCQ�����p8���   �QHP�ҋu���p8�H�QV�ҡp8�H�QVW�ҡp8���   ��U�R�Ѓ�$�M��}���_��^��]������U��p8�H��p  ��$�҅�u��]�Vh#���M������p8�P�E�R4Ph#���M���j �E�P�M�hicMCQ������p8���   �Q8P�ҋ�p8���   ��U�R�Ѓ��M�������^��]���������������U��p8�H��p  ��$�҅�u��]�Vhs���M��d����p8�P�E�R4Phs���M���j �E�P�M�hicMCQ�W����p8���   �Q8P�ҋ�p8���   ��U�R�Ѓ��M��E�����^��]���������������U��p8�H���  ]��������������U��p8�H��@  ]��������������U��p8�H���  ]��������������U��V�u���t�p8�QP��D  �Ѓ��    ^]������U��p8�H��H  ]��������������U��p8�H��L  ]��������������U��p8�H��P  ]��������������U��p8�H��T  ]��������������U��p8�H��X  ]��������������U��p8�H��\  ]�������������̡p8�H��d  ��U��p8�H��h  ]��������������U��p8�H��l  ]�������������̡p8�H���  ��U��p8�H�U���  ��VR�E�P�ыu��P���3����M��K�����^��]�����U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�H��$  ]��������������U��p8�H��(  ]��������������U��p8�H��,  ]�������������̡p8�H��0  ��p8�H��<  ��U��p8�H���  ]�������������̡p8�H���  ��U��p8�H���  ]������������������������������U��p8�H��  ]�������������̡p8�H��P  ��p8���   ���   ��Q��Y��������U��p8�H�A�U��� R�Ћp8�Q�Jj j��E�h��P�ыUR�E�P�M�Q�~���p8�B�P�M�Q�ҡp8�H�A�U�R�Ћp8�Q�J�E�P�у�,��]��V������F    �p8�H4���   �҉F��^����������V��V����p8�H4���   R��3����F�F^�������� �������������U����UR�UR�UR�UR�UR3��U��E��E���@R�U�R��3��}�gnol��H#E���]� ���������U��p8�P4�E�I���   P�EP�EP�EP�EP�EPQ�҃�]� ���������̡p8�P4�A���   P��Y����������̡p8�P4�A���   P��Y�����������U��p8�P4�E�I���   P�EP�EPQ�҃�]� ������U��p8�P4�E�I���   P�EPQ�҃�]� ����������U��p8�P4�E�I���   P�EP�EPQ�҃�]� ������U��p8�P4�E�I���   PQ�҃�]� �������������̡p8�P4�A���   P�у����������U��M��t#�U$��@R�U R�UR�UR�UR�UR�UR��]��U��E�@�p8�R4V�uQh�VP�A���   P�у�^]� ��������������V������F    �p8�H4���   �҉F����p8�Q4P���   �Ћp8�Q4���   ���ЉF��^�����������V��V����p8�H4���   R��3����F�F^�������U��p8�P4�E�I���   P�EPQ�҃�]� ����������U��p8�P4�E�I���   P�EPQ�҃�]� ����������U��p8�P4�E�I���   P�EPQ�҃�]� ���������̡p8�P4�A���   P�у����������U��p8�P4�E�I���   P�EP�EPQ�҃�]� ������U��p8�P4�E�I���   PQ�҃�]� ��������������� �������������U��p8�P4�E�I���   PQ�҃�]� ��������������U��p8�P4�E�I���   PQ�҃�]� ��������������U��p8�P4�E�I���   P�EPQ�҃�]� ����������U��p8�P4�E�I���   PQ�҃�]� ��������������U��p8�P4�E�I���   P�EPQ�҃�]� ����������U��V��V����p8�H4���   R��3����E�F�Ft	V���������^]� ���������������U���V�u�W�}�����Dz�F�_����D{:�F����$�@ �G��$�]��@ �E���������D{_�   ^��]�_3�^��]���������U���VW�M��0����E�}��t-�p8�Q4P�B�Ѓ��M��u�h���_3�^��]Ë�R(��p8�H0�QW�҃��M��tԋ�R Q�MQ���ҋ�p8�P�B �M��Ѓ��t�p8�Q0�Jx�E�PW�у��M������_��^��]�������U��p8�P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   �p8�Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� �p8�Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� �A���_3�^]� =cnys����_3�^]� ������V������p8�H0�Vh���҉F���F    ��^�����V��F�����t�p8�Q0P�B�Ѓ��F    ^�����̡p8�P0�A���   P�у����������U��p8�P0�E�I���   PQ�҃�]� �������������̡p8�I�P0���   Q�Ѓ���������̡p8�P0�A���   j j j j j j j j j4P�у�(������̡p8�P0�A���   j j j j j j j j j;P�у�(�������U��p8�P0�E�IPQ���   �у�]� ��������������U����E V��P�M������p8�E�Q�R4Ph8kds�M��ҡp8�E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M��Ȭ����^��]� ��������������̡p8�I�P0���   Q�Ѓ����������U��V��F��u^]� �p8�Q0�M ���   j j j j j Q�Mj QjP�ҡp8�H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uËp8�Q0P�B�Ѓ������̋A��u� �p8�Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5p8�v0Q�MQP���   R�U�R�Ћu�    �F    �p8���   j P�BV�Ћp8���   �
�E�P�у�$��^��]� �������U��p8�P0�E�I�RPQ�҃�]� �U��A��t)�p8�Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5p8�v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5p8�v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5p8�v0Q�MQPR�V\�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ�p8�P4�A�JhWVP�ы�ډ����ى_^]� �����U��A��u]� �p8�Q4�M�RhQ�MQP�҃�]� ����U��A��u]� �p8�Q4�M�RpQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ�p8�P4�A�JpWVP�ы�ډ����ى_^]� �����U���$VW��htniv�M��٨���p8�P�E�R4Phulav�M��ҡp8�P�B4hgnlfhtmrf�M��Ћp8�E�Q�R4Phinim�M��ҡp8�P�E�R4Phixam�M��ҡp8�P�E�R4Phpets�M��ҡp8�P�E�R4Phsirt�M��ҋE �}$=  �u�����t.�p8�QP�B4h2nim�M��Ћp8�Q�B4Wh2xam�M��ЋU�M�QR�E�P���K����p8���   P�B8�Ћp8���   �
���E�P�у��M������_��^��]�  ��������������U���$V��htlfv�M�芧���E�p8�P�B,���$hulav�M��Ћp8�E,�Q�R4Phtmrf�M����E�p8�P�B,���$hinim�M����E�p8�Q�B,���$hixam�M����E$�p8�Q�B,���$hpets�M��Ћp8�ED�Q�R4Phsirt�M��������E0��������Dzw���]8����Dzm�؋p8�E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R��������p8���   P�B8�Ћp8���   �
���E�P�у��M�蜦����^��]�@ �١p8�P�B,���$h2nim�M����E8�p8�Q�B,���$h2xam�M����V�����U���$V��hgnrs�M�������E�p8�E��E�   �Q���   �E�Pj�M��ҡp8���   ��U�R�ЋM�p8�M����E�   �B���   �M�Qj�M��ҡp8���   ��U�R�ЋU���M�QR�E�P��������p8���   P�B8�Ћp8���   �
���E�P�у��M��z�����^��]� �U���$V��hCITb�M������p8�P�E�R8PhCITb�M��ҡp8�P�E�R4Phsirt�M��ҡp8�P�E�R4Phulav�M��ҋM�E�PQ�U�R�������p8���   P�B8�Ћp8���   �
���E�P�у��M��ɤ����^��]� U��E��Vj ��P�M�Q�M�e����UPR���)�����p8�H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�O���]�( �����������U��E,��Pj ���T$�U�$hrgdf�E$�� �������������\$�E�����\$�M���\$�E�$R�����]�( ���U��E,��Pj ���T$�U�$htcpf�E$�� ��������\$�E���\$�}�\$�E�$R����]�( ���������������U��Q��u3�]� �E�E�H� V�5p8�v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5p8�v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5p8�v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5p8�v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5p8�^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� �p8�[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=p8�0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5p8�v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3�W��u3��,�E�H� �5p8�v0Q�MQPR�V,��3Ƀ�9M������p8�M�B�P0VQ�M�ҋ�_^]� ����U��AV��u3��"�M�Q�	�5p8�v0R�URQP�F,�Ѓ����p8�Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A��V��u3��"�M�Q�	�5p8�v0R�U�RQP�F0�Ѓ����p8�E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U��V�U��]�W��t$�E�H� �=p8�0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=p8�0Q�M�QPR�W0�҃���tˋV��tċE�H� �5p8�v0Q�M�QPR�V0�҃���t��p8�P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A�U�V�U�W�]���u3��&�M�Q�	�5p8�v0R�U�R�U�RQP�F<�Ѓ����E�}���t�p8�Q�RH�M�QP���ҋE���t�p8�E��Q���$P�B,����_��^��]� U��p8�P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR���o���^]�  ����������U��p8��P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�K���^]�< ������U��p8��P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P�����^]�$ �����������U��p8��P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P�C���^]�$ ��������������U��p8��P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� ����������\$�E���\$�}�\$�$P����^]�$ ���������������U��p8�� V��H�A�U�R�ЋM�E��Qj �U�RP�M�Q�M��B���UPR��������p8�H�A�U�R�Ћp8�Q�J�E�P�у���^��]� ������������U���dV��M��Oz���p8�Q���   P�EP�M�Q�M��P�M���z���M��{��j j �E�P�M���{���MPQ�������p8���B�P�M�Q�҃��M���z���M���z����^��]� �����U���P��EV�]���W�}����t�p8�Q���$P���   �����]���p8�U��UЍE��]ȋQ�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F�U��u_^��]� �M�E�Q�	�5p8�v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E�M���u�p8�H���   �҅�u��]� SVW���L�����htlfv�MЉu�Z����E�}�p8�X�U�����$�<* �]��G�$�.* �}�S,�M��$hulav�ҡp8�P�B4hmrffhtmrf�M��Ћ}��p8�M�Y���$��) �]��G�$��) �}�S,�M��$hinim�ҋ}��p8�M�X���$�) �]��G�$�) �}�S,�M��$hixam����p8�P�B,���$hpets�M��Ћp8�Q�B4j hdauq�M��Ћp8�Q�B4Vhspff�M��Ћp8�E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R�n����p8���   P�B8�Ћp8���   �
���E�P�у��M�����_��^[��]� U��E��V���u�p8�H���   �҅�u^��]� ���~����E�F��u3��"�M�Q�	�5p8�v0R�U�RQP�F0�Ѓ����E������M������\$�M��$謷  ��M��P�Q�P�Q�@�A��^��]� ����������U���0��p8�]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP�����p8�Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5p8�v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� �p8�Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� �p8�Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U��p8�P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� �p8�Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5p8�v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M����  �MQ�U�R�M��H�  ��tm�}��E��tN�p8���   P�BH�ЋM��I����tQ�W�7�p8�[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M��۴  ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5p8�v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� �p8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �p8�Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� �p8�Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uËp8�Q0P�BX�Ѓ�������U��A��u]� �p8�Q0�M�RLQ�MQP�҃�]� ����U��A��u]� �p8�Q0�M�RP��   �QP�҃�]� ��U��A��u]� �p8�Q0�M�RPQP�҃�]� ��������U��A��u]� �p8�Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U��p8V�u�VW���H4�R�ЋE�F    �~�H� �p8�R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� �p8�Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I�p8�R0P�EPQ���   �у�]� ������̡p8�I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u�`8� �p8�R0�I�R@V�uVP�EPQ�҃�^]� �����������U��p8�P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U��p8�P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5p8�v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� �p8�R0j j j j j j j P�A���   jP�у�(]� �����������U��E� �p8�R0j j j j j jj P�A���   jP�у�(]� �����������U��E� �p8�R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� �p8�R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R諈���M�蓈����^��]� ����������U��E�P� V�5p8�v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5p8�v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5p8�v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5p8�v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U��p8�P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U��p8�UVj j j j j R��H0�E�Vj P���   jR�Ћp8�Q0�E�N�RtPQ�҃�0^]� ��U��p8�P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡p8�P0�A���   j j j j j j j j jP�у�(�������U��p8�P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡p8�P0�A���   j j j j j j j j j(P�у�(�������U��p8�P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U��p8�P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡p8�P0�A���   j j j j j j j j jP�у�(������̡p8�P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���t�p8�P���   j j���Љ�u��t�p8�Q���   j j���Љ�p8�Q0�E��H�R`VWQ�҃�_^[��]� �U��p8�P0�E�I���   P�EP�EPQ�҃�]� �����̡p8�P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V������p8�H0�Vh���҉F3��F�F������F   ��^�������V��F�����t�p8�Q0P�B�Ѓ��F    ^������U��E�UVj ��MP�EQ3�9MR��Pj �F    ��
Q��������t�~ t
�   ^]� 3�^]� �U��E�A�I��u3�]� �p8�B0Q�H�у�]� ����U��p8�P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   �p8�Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tK��B����^[]� �~ t6��������t+�F    ^�   []� =atnit�MQS���/���^[]� ^3�[]� �U��V��~ ��   W�}����   �$�8��E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN�p8�M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W訷�����F    _^]� d�r�������������������U��V��~ �  �E W�}�E����   �$������]������   �   ���]����A��   �   ���]����A��   �r���]������   �`�E������A��uN��������   �C�E��������u1������A{{�*�E���������E������A�����]����DzU����ءp8�U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W�S������F    _^]�$ �I ��������������&�������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� ��H�H�H�������������VW��3���9~u�p8�H4�V�R�Ѓ��~�~_^����U��p8�P4�E�I�RtPQ�҃�]� �U��U��t3�A�p8�I0R���   P�ҋp8�Q0�M���   QP�҃�]� �p8�P0�E�I�R|PQ�҃�]� ������̡p8�P4�A�JP�у������������̡p8�P4�A�JP�у������������̡p8�P4�A�JP�у������������̡p8�P4�A�J|P�у������������̡p8�P4�A���   P�у����������U��p8�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U��p8�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U��p8�P4�E�I�R PQ�҃�]� �U��p8�P4�E�I�R$PQ�҃�]� �U��p8�P0�E�I���   P�EP�EP�EPQ�҃�]� ��U��p8�P4�E�I���   PQ�҃�]� ��������������U��p8�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��p8�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��p8�P4�E�I�R(PQ�҃�]� �U��p8�P4�E�I�R,P�EP�EPQ�҃�]� ���������U��p8�P4�E�I�R0P�EPQ�҃�]� ������������̡p8�P4�A�J4P��Y��������������U����UV��EP�M�Q�NR�E�    �E�    �����p8�H4�V�AR�Ћp8�Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃� �} ^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ��������������U��p8�P4�E�I�R8PQ�҃�]� �U��p8�P4�E�I�R<PQ�҃�]� �U��p8�P4�E�I���   P�EPQ�҃�]� ���������̡p8�P4�A�J@P�у�������������U��p8�P4�E�I�RDP�EPQ�҃�]� �������������U��p8�P4�E�I�RHP�EPQ�҃�]� �������������U��p8�P4�E�I�RLP�EPQ�҃�]� �������������U��p8�P4�E�I�RPP�EPQ�҃�]� �������������U��p8SV�uW�����   �QV�҃�����   �p8���   �]�QS�҃�S��uA�p8���   �Q@�ҋءp8���   �Q@V�ҋp8�Q4�JPSP�GP�у�_^[]� �p8���   �H�у���uD�p8���   �H8S�ыp8�؋��   �H@V�ыp8�J4�WSP�AHR�Ѓ�_^[]� h@�h}  ��   �p8���   �BV�Ѓ�����   �p8���   �]�BS�Ѓ�S��uC�p8���   �B@�Ћp8���   �؋B8V�Ћp8�Q4�JLSP�GP�у�_^[]� �p8���   �H�у���uD�p8���   �H8S�ыp8�؋��   �H8V�ыp8�J4�WSP�ADR�Ѓ�_^[]� h@�h�  �
h@�h�  �p8�Q��0  �Ѓ�_^[]� �U��p8�P4�E�I��  P�EP�EP�EPQ�҃�]� ��U��p8�P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U��p8�P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡p8�P4�A�J`P��Y�������������̡p8�P4�A�JdP�у�������������U��p8�P4�E�I��   P�EP�EP�EPQ�҃�]� ��U��p8�P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U��p8�P4�E�I�RhP�EPQ�҃�]� �������������U��V�uW��t��؉�}��t��ډ�p8�P4�A�JhWVP�у���t��ډ��t��ى_^]� �U��V�uW��t��؉�}��t��ډ�p8�P4�A�JpWVP�у���t��ډ��t��ى_^]� �U��p8�P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   �p8�V�H4�AR�Ѓ} t �p8�Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �Lt��P�M�Q�N�U�R�����p8���   ��U�R�Ѓ��M��]t��^��]� ������U��p8�P4�E�I�RlPQ�҃��   ]� ������������U��p8�E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U��p8�P4�E�I���   P�EP�EPQ�҃�]� �����̡p8�P4�A���   P�у���������̸   ����������̸   �����������U��p8V��H4�V�A$h�  R�Ћp8�Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U��p8�P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U��p8�P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���t�p8�P���   j j���Љ�u��t�p8�Q���   j j���Љ�p8�Q4�E��H�RpVWQ�҃�_^[��]� �U��Q�p8�P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t�p8�U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  �p8�Q���   j j���Ћp8�Qj �؋��   j���Ћp8�Qj �E����   j���Ћp8�Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���Y���P���1���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� �p8�Q���   j hIicM���ЋWP�B ����_^[��]� �������������U��p8�P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��*o���p8�Q4�JlP�FP�у��M��Lo��^��]��������V������p8�H0�Vh���҉F���F    ����F   ��^��������V��F�����t�p8�Q0P�B�Ѓ��F    ^������U��p8�P�B VW�}�����=cksat`=ckhct�MQW��譾��_^]� �Nj j j j j j �F   �p8�B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U��p8�H���  ]��������������U��p8�H0���   ]��������������U��p8�H0�U�E��VWRP���   �U�R�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�_��^��]������������U��p8�H0���   ]��������������U��p8�H0���   ]��������������U��Ej0P貞����]��������������U��Ej0P�;����P艞����]�����U��E�M��j0PQ�U�R�;����P�^����p8�H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P��<����P�����p8�Q�J�E�P�у���]��U��Ej$P����3Ƀ�������]����U��Ej$P��:����P�ɝ��3Ƀ�������]�����������U��E�M��Vj$PQ�U�R��:����P荝���p83Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P��;����P�9����p83Ƀ��B�P����M�Q�҃���^��]����U��p8�H�U�E���   RPj �у�]���������������U��p8�H�U�ER�UP���   Rj �Ѓ�]�����������U��p8�P4�E�I�R,P�EP�EPQ�҃�]� ���������U��p8�P4�E�I�R0P�EPQ�҃�]� ������������̡p8�P4�A�J4P��Y��������������U��U��V��EP�M�QR���d����p8�H0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ��} ^t(�} t(�E�M�;�~<�U��;�}3�E�M�;�~)�U���} u�E�M�;�~�U��;�}�   ��]� 3���]� �����������U��ESVW�؅�u�Y�p8�P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� �p8�Q���   j hIicM����;�u�p8�Q���   j h1icM���Шu��3_^�   []� �����U��p8�P�BT��(V�uhfnic���Ѕ�t�p8�Q�ȋ��   j
�Ѕ���   �p8�Q�RPhfnic�E�P����P�M���h���M��i���u�E�P���	i���M���h���p8�Q�B ���Ѓ��t�p8�Q�B ���Ѕ�u�p8�Q�B$hfnic���Ћp8�E�Q�R8Pj
����^��]���������U��p8�P0�E�IP�EP�EP�EPQ���   �у�]� ��U��p8�P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U��p8�P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡p8�I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V������p8�H0�WVh���ҋ}�F�E�F    �F   ����F�p8�Q���   ��j hmyal���ЉF��t��t�F    �p8�Q���   j
hhfed���ЉF_��^]� �����������U��p8�P�B VW�}�����=ytsdt�MQW������_^]� �p8�B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸ ������������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&�p8�R0j j j j j j P���   j jQ�Ѓ�(�p8�Q�J�E�P�ыp8�B�P�M�Q�ҋF����t �p8�Q0�RHj �M�Qj jj?j P�҃��p8�H�A�U�WR�Ћp8�Q�J�E�P�ыF����u3��;�p8�E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(�p8�Q�J�E�P�у���_u3�^��]Ëp8�B�P�M�Q�ҋF����t �p8�Q0�RHj �M�Qj j j8j P�҃��p8�H�A�U�R�ЋF����t�p8�Q0jP�BP�Ѓ��p8�Q�J�E�P�у��M��c��Ph   h  K j;�U�Rh	��h�  ��跶���p8�H�A�U�R�Ѓ��M���c���F��t�p8�Q0P�BX�Ѓ��F��t�p8�Q0P�BX�Ѓ��F��t'�p8�Q0j j j j j jj j jP���   �Ѓ�(j�v$葔�����   ^��]�����U���SV��W�~j����e����V�^(3ۉ^4�^8�^<�p8�H0�Ah�   R�Ћp8�Q�J�E�P�ыp8�B�PSj��M�h�Q�҃�SS�E�P�M�Q���E��  �]��i����p8�B�P�M�Q�҃�Sj���
e��_^[��]���̍A�������������U��VW��~4 tA�I �p8�H��0  h@�hj  ��j
�o����p8�HP�V �AR�Ѓ���uQ9F4up8�QP�Bh�~0���Ѓ~4 t;�p8�Q��0  h@�h�  �Ћp8�QP�Bl�������m���_3�^]� �M�U�N8�V4�p8�PP�Bl�~0���Ѓ~4 t%j
�Ӝ���p8�QP�F �JP�у���u�9F4uۋp8�BP�PhS���ҋ^<�F<    �p8�PP�Bl���Ћ�[_^]� ��U��p8�P�B ��@VW�}�����=MicMtI=fnic��   j�M��a���uP���Ma���M��5a���p8�Q�B4jj����_�   ^��]� �p8�Q���   j hIicM����=�����   htats�M��`���p8�Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    �̴���p8���   �
�E�P�у��M��`���F�F   ��t�p8�J0�QP�҃��EPW���a���_^��]� ���������U��E��V��t3�^]� j�N�b��j�J����F    �v����t�p8�H0�QV�҃��   ^]� ��������������j���fb��j�������3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�u���]� �U��Q�Q��u3���]� �E�H� V�5p8Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9�p8�Q�M�RQP�ҋE�����t�p8�QW��P�B��W��g����_��^��]� ������U��p8��V��H�A�U�R�ЋU���M�QR���D�������u�p8�H�A�U�R�Ѓ�3�^��]� �M�Q�M��>���p8�B�P�M�Q�҃���^��]� �������U��p8��V��H�A�U�R�ЋU���M�QR��������M��p8�P�R8�E�PQ�M�ҡp8�H�A�U�R�Ѓ���^��]� �������������U���V��M��<���M�E�PQ��������p8���B�U�@<�M�Q�MR�ЍM���<����^��]� ����U��p8�P�E���   Vj ��MP��h���h  �j j jj P�EP���c���^]� ��������������U��p8V�uW�����   �QV�҃�V��u,�p8���   �Q@�ҋp8�Q4�J P�GP�у�_^]� �p8���   �H�у���u.�p8���   �H8V�ыp8�J4�WP�A$R�Ѓ�_^]� �p8�Q��0  h@�h	  �Ѓ�_^]� �����U���4�p8�H�QSVW�}W�ҡp8�P�u���   ��3�SS�Ή]�Ћp8�QS�E����   j���Ћ�;��L  �d$ �} ~l�p8�Q�J�E�P�ыp8�B�Pj j��M�h�Q�ҡp8�P�B<�����Ћp8�Q�RLj�j��M�QP���ҡp8�H�A�U�R�Ѓ��p8�Q0�E����   VP�M�Q�ҋ�p8�H�A�U�R�Ћp8�Q�J�E�PV�ыp8�B�P�M�Q�ҡp8�P�B<�����Ћp8�Q�RLj�j��M�QP���ҡp8�H�A�U�R�Ћp8�Q�u���   �E��j ��
S���Ћp8�Q���   �E�j �CP���ҋ����������_^[��]����������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR��荱��^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�O���^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P�B���]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P����]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P�j���]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� ��������\$�E���\$�}�\$�$P�K���]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�_���^]� ����������U��Q��u3�]� �E�E�H� V�5p8�v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U��p8�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U��p8�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U��p8��P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�^����D{�   ^]� ��^]� ������U���0��p8�U�V�U���M�]�P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A����  ^��]� ��������U��� ��p8�]�V���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�@�Q�A����  ^��]� �����U���VW�}�M�;}us�p8�P�u���   j htsem���Ѕ�uS�p8�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��'�����t�E�M�P�w  _�   ^��]� _3�^��]� U���VW�}�M�;}us�p8�P�u���   j htsem���Ѕ�uS�p8�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�������t�E�M�P��  _�   ^��]� _3�^��]� U���SVW�}��;}uz�p8�P�u���   j htsem���Ѕ�uZ�p8�QP���   hrdem���Ѕ�u=��M�Q�]��M�U�R�}��E�蕲����t�E������$�  _^�   [��]� _^3�[��]� ��������U���4�ESW�}�M�;�t;Et	;E��   �p8�P�]���   j htsem���Ѕ���   �p8�QP���   hrdem���Ѕ�uj�M��U�U܉E��UԉE��]̉E�M�E�P�M�Q�M�U�U�R�E�P�}�������t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�}��;}��   �p8�P�u���   j htsem���Ѕ�uj�p8�QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}��x�����t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h���� ������������������U��p8��0VW���H�A�U�R�Ћp8�Q�J�E�P�ыE���U�RP�M�Q�M�<����p8�J�U�RP�A�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�ҡp8�H�Q��V�ҡp8�H�A�U�VR�Ѓ�����  �p8�Q�J�E�P�у�_^��]� ������������U���SVW�}��;}��   �p8�P�u���   j htsem���Ѕ�ue�p8�QP���   hrdem���Ѕ�uH�p8�Q�J�E�P�ыM���U�R�E�P�}��E�    �-�����u �p8�Q�J�E�P�у�3�_^[��]� ���U��R�������  �p8�H�A�U�R�Ѓ�_^�   [��]� ��U��V�u���  ��^]� �����������U���L�p8SV��H�A�U�R�Ћp8�Q�J3�Sj��E�h�P���F(�����S�U�SR�E��  �]����  P�E�P�n�����P�M�Q�1����P�U�R���b����p8�H�A�U�R�Ћp8�Q�J�E�P�ыp8�B�P�M�Q�҃�htats�M��MP���p8�P�B0jj�M����F(�p8�Q�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]��`����p8���   �
�E�P�у�9^4t^�p8�BP�PhW�~0���ҋF4;�t�N8Q�Ѓ��F<�^8�^4��p8�B��0  h@�h�  �у��p8�BP�Pl����_�M��O��^[��]� ������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�E�Y����D{�   ]� �����������U�����u�E�    �Y�E�Y�E�Y]� ��u-�E�Y����Dz�E�Y����Dz�E�Y����D{�   ]� �����U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR菝������t�   ^]� �������������U��V��~ ��u�p8�H4�V�R�Ѓ��E�F    �F    t	V�W������^]� �������U��V��F�����t�p8�Q0P�B�Ѓ��E�F    t	V��V������^]� ��������������U���V��3ɍF��H������p8�M��M����   �RQ�M�QP�ҡp8���   ��U�R�Ѓ���^��]��������������U��V�����u �    �p8�H�A���UVR�Ѓ��#��u�p8�Q�Rx�EP�N�҅�t�   �p8�H�A�UR�Ѓ�^]� �������hx8PhD ��u  ���������������U��Vhx8h�   hD ���u  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vhx8h�   hD ���Vu  ����t���   ��t�M�UQR����^]� 3�^]� �������������U���VWhx8h�   hD ���u  ��3���;�tH9��   t@�M�E�E��E�E��E�E��E�PQ�0�  ����t�UR���   �E�P����_^��]� _3�^��]� �����U��Vhx8h�   hD ���t  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vhx8h�   hD ���6t  ����t���   ��t�MQ����^]� ��������U��Vhx8h�   hD ����s  ����t���   ��t�MQ����^]� ��������U��Vhx8h�   hD ���s  ����t���   ��t�MQ����^]� ��������U��Vhx8h�   hD ���vs  ����t���   ��t�MQ����^]� ��������h|8PhD �@s  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h|8jhD �lr  ����t
�@��t]��3�]��������Vh|8j\hD ���<r  ����t�@\��tV�Ѓ���^�����Vh|8j`hD ���r  ����t�@`��tV�Ѓ�^�������U��Vh|8jdhD ����q  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh|8jhhD ���q  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh|8jlhD ���\q  ����t�@l��tV�Ѓ�^�������U��Vh|8h�   hD ���&q  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh|8h�   hD ����p  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh|8jphD ���p  ����t�@p��t�MQV�Ѓ�^]� ��8^]� ��U��Vh|8jxhD ���Ip  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh|8jxhD ���	p  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh|8jxhD ����o  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h|8jhD �oo  ����t	�@��t��3��������������U��V�u�> t+h|8jhD �3o  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h|8jhD ��n  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh|8jhD ���n  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh|8jhD ���in  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh|8j hD ���,n  ����t�@ ��tV�Ѓ�^�3�^���Vh|8j$hD ����m  ����t�@$��tV�Ѓ�^�3�^���U��Vh|8j(hD ����m  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh|8j,hD ���ym  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh|8j(hD ���9m  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh|8j4hD ����l  ����t�@4��tV�Ѓ�^�3�^���U��Vh|8j8hD ���l  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh|8j<hD ���il  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh|8jDhD ���,l  ����t�@D��tV�Ѓ�^�3�^���U��Vh|8jHhD ����k  ����t�M�PHQV�҃�^]� U��Vh|8jLhD ����k  ����u^]� �M�PLQV�҃�^]� �����������U��Vh|8jPhD ���k  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh|8jThD ���Lk  ����u^Ë@TV�Ѓ�^���������U��Vh|8jXhD ���k  ����t�M�PXQV�҃�^]� U��Vh|8h�   hD ����j  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh|8h�   hD ���j  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh|8h�   hD ���Fj  ����u^]� �M���   QV�҃�^]� �����U��Vh|8h�   hD ���j  ����u^]� �M���   QV�҃�^]� �����U��Vh|8h�   hD ����i  ����u^]� �M���   QV�҃�^]� �����U��Vh|8h�   hD ���i  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh|8h�   hD �Ei  ����u�p8�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћp8�Q�u���BV�Ћp8�Q�BVW�Ћp8�Q�J�E�P�у�_��^��]��U��Vh|8h�   hD ���h  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh|8h�   hD ���fh  ����t���   ��t�MQ����^]� 3�^]� �U��Vh|8h�   hD ���&h  ����t���   ��t�MQ����^]� 3�^]� �U��Vh|8h�   hD ����g  ����t���   ��t�MQ����^]� 3�^]� �Vh|8h�   hD ���g  ����t���   ��t��^��3�^����������������U��Vh|8h�   hD ���fg  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh|8h�   hD ���g  ����t���   ��t�MQ����^]� ��������U��Vh|8h�   hD ����f  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh|8h�   hD ���f  ����t���   ��t��^��3�^����������������VW��3����$    �h|8jphD �?f  ����t�@p��t	VW�Ѓ����8�8 tF��_��^�������U��SW��3�V��    h|8jphD ��e  ����t�@p��t	WS�Ѓ����8�8 tqh|8jphD �e  ����t�@p��t�MWQ�Ѓ������8h|8jphD �e  ����t�@p��t	WS�Ѓ����8V���7�����tG�]����E^��t�8��~=h|8jphD �>e  ����t�@p��t	WS�Ѓ����8�8 u_�   []� _3�[]� ����������U��Vh|8j\hD ����d  ����t3�@\��t,V��h|8jxhD ��d  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh|8j\hD ���d  ����t3�@\��t,V��h|8jdhD �gd  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh|8j\hD ���&d  ����tG�@\��t@V�ЋEh|8jdhD �E��E�    �E�    ��c  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh|8j\hD ���c  ����t\�@\��tUV��h|8jdhD �c  ����t�@d��t
�MQV�Ѓ�h|8jhhD �^c  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh|8j\hD ���c  ������   �@\��t~V��h|8jdhD ��b  ����t�@d��t
�MQV�Ѓ�h|8jhhD ��b  ����t�@h��t
�URV�Ѓ�h|8jhhD �b  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh|8jthD ���fb  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h|8j`hD �.b  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�8���_�����^��]� ������U���Vh|8h�   hD ����a  ����tR���   ��tH�MQ�U�R���ЋuP������h|8j`hD �a  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�BQ�Ѓ����������������U��p8�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U��p8�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��p8�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��p8�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U��p8�PX�EPQ�J�у�]� ����U��p8�PX�EPQ�J�у�]� ����U��p8�PX�EPQ�J�у�]� ����U��p8�PX�EPQ�J�у�]� ����U��p8�PX�EPQ�J$�у�]� ����U��p8�PX�EPQ�J �у�]� ����U��p8�PD�EP�EPQ�J�у�]� U��p8�HD�U�j R�Ѓ�]�������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�HD�	]��U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�HD�U�j R�Ѓ�]�������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�U�HD�Rh2  �Ѓ�]����U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�U�HD�RhO  �Ѓ�]����U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�U�HD�Rh'  �Ѓ�]����U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�HD�j h�  �҃�����������U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�HD�j h:  �҃�����������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E��p8���   �R�E�Pj�����#E���]�̡p8�HD�j h�F �҃�����������U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�HD�j h�_ �҃�����������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E��p8�E�    ���   �R�E�Pj������؋�]� ̡p8�PD�B$Q�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ���������������̡p8�PD�B(Q�Ѓ���������������̡p8�PD�BQ�Ѓ����������������U��p8�E�PH�B���$Q�Ѓ�]� ���������������U��p8�PH�EPQ���   �у�]� �U��p8�PH�EPQ���  �у�]� �U��p8�PH�EPQ���  �у�]� �U��p8�PH�EP�EPQ��  �у�]� �������������U��p8�PH�EP�EPQ��  �у�]� ������������̡p8�PH���  Q�Ѓ�������������U��p8�PH�EPQ���  �у�]� ̡p8�PH���   j Q�Ѓ�����������U��p8�PH�EPj Q���   �у�]� ��������������̡p8�PH���   jQ�Ѓ�����������U��p8�PH�EPjQ���   �у�]� ��������������̡p8�PH���   jQ�Ѓ����������U��p8�PH�EPjQ���   �у�]� ���������������U��p8�PH�EP�EPQ���   �у�]� �������������U��p8�PH�EP�EPQ���   �у�]� ������������̡p8�PH���   Q�Ѓ�������������U��p8�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���@���������t�E�p8�QH���   PVW�у���_^]� �����U��EVW���MPQ�L���������t�M�p8�BH���   QVW�҃���_^]� ̡p8�PH���   Q�Ѓ������������̡p8�PH���   Q�Ѓ�������������U��p8�PH�EPQ���   �у�]� �U��p8�PH�EPQ���   �у�]� �U��p8�PH�EP�EPQ��8  �у�]� �������������U��p8�PH�EP�EPQ��   �у�]� ������������̡p8�PH���  Q�Ѓ������������̡p8�PH���  Q�Ѓ������������̡p8�PH���  Q�Ѓ������������̡p8�PH��  Q�Ѓ������������̡p8�PH��  Q�Ѓ�������������U��p8�PH�EP�EPQ��  �у�]� �������������U��p8�PH�EP�EP�EPQ��   �у�]� ���������U��p8�PH�EP�EP�EP�EPQ��|  �у�]� �����U��p8�PH�EPQ��  �у�]� ̡p8�PH��T  Q�Ѓ�������������U��p8�PH�EP�EPQ��  �у�]� �������������U��p8�PH�EPQ��8  �у�]� �U��p8�PH�EPQ��<  �у�]� �U��p8�PH�EPQ��@  �у�]� �U��p8�PH�EP�EP�EPQ��D  �у�]� ��������̡p8�PH��L  Q��Y��������������U��p8�PH�EPQ��H  �у�]� ̡p8V��H@�Q,WV�ҋp8�Q��j �ȋ��   h�  �Ћp8�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡p8�P@�B,Q�Ћp8�Q��j �ȋ��   h�  �������U��p8�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��p8�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��p8�PH�EP�EP�EPQ��   �у�]� ��������̡p8�HH��  ��U��p8�HH��  ]��������������U��p8�E�PH��$  ���$Q�Ѓ�]� �����������̡p8�PH��(  Q�Ѓ�������������U��p8�PH�EP�EPQ��,  �у�]� �������������U��p8�E�PH�EP�E���$PQ��0  �у�]� ���̡p8�PH���  Q�Ѓ������������̡p8�PH��4  Q�Ѓ������������̋��     �������̡p8�PH���|  jP�у���������U��p8�UV��HH��x  R��3Ƀ������^��]� ��̡p8�PH���|  j P�у��������̡p8�PH��P  Q�Ѓ������������̡p8�PH��T  Q�Ѓ������������̡p8�PH��X  Q�Ѓ�������������U��p8�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡p8�PH��`  Q�Ѓ�������������U��p8�PH�EPQ��d  �у�]� �U��p8�E�PH��h  ���$Q�Ѓ�]� ������������U��p8�E�PH��t  ���$Q�Ѓ�]� ������������U��p8�E�PH��l  ���$Q�Ѓ�]� ������������U��p8�PH�EPQ��p  �у�]� �U��p8�PH�EP�EP�EP�EPQ���  �у�]� �����U��p8�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U��p8�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E�p8�HH�E���   R�U���$P�ERP�у�]����������������U���E�M� �謴  �M;�|�M;�~��]�����������U��p8�PH�E���   Q�MPQ�҃�]� ������������̡p8�PH���   Q��Y�������������̡p8�PH���   Q�Ѓ������������̡p8�PH���   Q��Y��������������U��p8�PH�EP�EPQ���   �у�]� �������������U��p8�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡p8�PH��t  Q��Y�������������̋�� ,��@    ��,��p8�Pl�A�JP��Y��������U��p8V��Hl�V�AR�ЋE����u
�   ^]� �p8�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uËp8�QlP�B�Ѓ�������U��p8�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E�p8�HH�ER�U���$P���  R�Ѓ�]����U��p8�HH���  ]��������������U��p8�HH���  ]��������������U��U0�E(�p8�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U��p8�HH���  ]��������������U��p8�E�PH�EP���$Q���  �у�]� ��������U���SV���&  �؉]����   �} ��   �p8�HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}���&  ����   �]��I �E�P�M�Q�MW�'  ��ta�u�;u�Y�I ������u�E�������L�;Ht-�p8�Bl�S�@����QR�ЋD������t	�M�P�c&  F;u�~��}��MG�}��.&  ;��v����]�_^��[��]� ^3�[��]� ��������������U����p8SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u�p8�HH���  �'��u�p8�HH���  ���ušp8�HH���  S�ҋȃ��E��t�W��%  �p8�HH���   h�  S3��҃����  ���_�u����    �p8�Hl�U�B�IWP�ы�������   �p8�F�J\�UP�A,R�Ѓ���t�K�Q�M�%  �p8�F�J\�UP�A,R�Ѓ���t�K�Q�M��$  �E��;Pt&�F�p8�Q\�J,P�EP�у���t	�MS�$  �p8�v�B\�M�P,VQ�҃���t�M�CP�$  �p8�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U��p8�HH���   ]�������������̡p8�PH���   Q��Y��������������U��p8�HH���  ]��������������U��p8��P���   V�uW�}���$V�����E������At���E������z����؋p8�Q�B,���$V����_^]����������������U���0��p8�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١p8�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U��p8�HH�]��U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�HH�h�  �҃�������������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�HH�Vh  �ҋ�������   �EPh�  ��������t]�p8�QHj P���   V�ЋMQh(  �V�������t3�p8�JH���   j PV�ҡp8���   �B��j j���Ћ�^]áp8�H@�QV�҃�3�^]�������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�HH�Vh�  �ҋ�����u^]áp8�HH�U�E��  RPV�у���u�p8�B@�HV�у�3���^]�������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�HH�I]�����������������U��p8�H@�AV�u�R�Ѓ��    ^]��������������U��p8�PH�EPQ���  �у�]� �U��p8�PH�EPQ���  �у�]� ̡p8�PH���  Q�Ѓ�������������U��p8�HH���  ]��������������U��p8�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡p8�PH���  Q�Ѓ�������������U��p8�PH�EP�EPQ���  �у�]� ������������̡p8�PH��  Q�Ѓ�������������U��p8�PH�EP�EP�EPQ���  �у�]� ��������̡p8�PH���  Q�Ѓ������������̡p8�PH���  Q�Ѓ�������������U��p8�PH�EPQ��  �у�]� �U��p8�PH�EPQ��  �у�]� ̋������������������������������̡p8�HH���  ��U��p8�HH���  ]��������������U��p8�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U��p8�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡p8�PH��,  Q�Ѓ�������������U��p8�PH�EPQ��X  �у�]� ̡p8�PH��\  Q�Ѓ�������������U��p8�HH��0  ]��������������U��p8��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �������������   �p8�HH���   j VW�҃��M��s���p8�P�E�R0Ph�  �M����E�p8�P�B,���$h�  �M��Ћp8�Q@�J(j �E�PV�у��M��|��^�   _��]� ^3�_��]� �����U��S�]�; VW��u7�p8�U�HH���   RW�Ѓ���u�p8�QH���   jW�Ѓ���t�   �����   �p8�QH���   W�Ѓ��} u(�p8�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;�p8�U�HH�ER�USP���  VRW�Ћp8���   �B(�����Ћ���uŃ; u�p8�QH���   W�Ѓ���t3���   �W��u1�p8�QH���   �Ћp8�E�QH���   PW�у�_^[]� �p8�BH���   �у��} u0�p8�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� �p8�QH�h  �Ћ؃���u_^[]� �p8���   �u�Bx���Ћp8���   P�B|���Ѕ�tU�p8�E�QH�MP�Ej Q���  VPW�у���t�p8���   �ȋBHS�Ћp8���   �B(���Ћ���u�_^��[]� ��������������U��EV���u�p8�HH���  �'��u�p8�HH���  ���u�p8�HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D�p8�HH���   S�]VWh�  S�ҋ�p8�HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��.
  �p8���   �B���Ћp8=�  ��  �QH���   Wh:  S�Ћp8�QH�E����   h�  S�Ћp8�QHW�����   h�  S�uԉ}��Ћp8�QH�E苂  S�Ћp8�QH�EЋ��  S�Ѓ�(�E��E�8���~~�M���M�I �MЅ�tMj�W�Au  ���t@�@�Ẽ|� �4�~����%�������;�u/���P~  ;E�~�E؋��~  E���E�;Pu�E���E��E�G;}�|��}� tv�u�j S�����������  ���������tV�������}�;�uK�p8�H���  �4�h@���h�  V�҃��E���N  �M�PVP����P�ׄ  ����}ܡp8�H���  �4�h@���h�  V�҃��E����  �M�3�;�t;�tVQP��  ���E�;�~-�p8�Qh@���h�  P���   �Ѓ��E�;���  �p8�E��QH��  j�PS�у�����  �u�;�tjS����������{  ��������E���}�p8�BH���   Wh�  S�у�3�9}ԉE�}��`  �}���}Ȑ�MЅ��R  �U�j�R�Js  ����>  �M̍@�|� ���]�~����%�������9E���  ���|  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����E؅��9  �+U�j��PR�M��5`  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$�4c�U����4�"�M����t��U����t�
�M����t�M���;]�|��E܃�F;]؉M��	����U�;U��
  �U�R����E�P�����M�Q������_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���P�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@��;EԉE��}�������U�R�����E�P�������  ���   �B����=  ��  �p8�QH���   j h(  S�Ћp8�QH�����   h(  S�ЋЃ�3��U؅�~'����    �ǅ�t�|� t�4N��tN�@;�|�u��u܋p8�Q���  �4v�h@���hK  V�Ѓ��E�����   �M��t��tVQP��  ���u؋p8�Q���  �h@���hP  V�Ѓ��E���tP��t��tVWP�֛  ���M����+p8�RH��PQ�E���   S�Ѓ���u�M�Q����U�R�����_^3�[��]áp8�HH���   j h�  S�҉E��p8�HH���   j h(  S��3�3���3�9]؉E��}ĉ]��7  �U��څ��  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�F@F����;�|��}ă|� ts�U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�F�v�Ћ��A�B�A�B�A�B�A�B�I�J�U�F<ډ}�C;]؉]�������M�3�3�;�~�U����$    ��t���   @;�|��U�R�������E�P�����_^�   [��]�]�]�]�]������������U��E� �M+]� ���������������U��V��V�,��p8�Hl�AR�Ѓ��Et	V�������^]� ���������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�p8���   P�B@��]� �E��t�p8���   P�BD��]� �p8���   R�PD��]� �����U��p8�P@�Rd]�����������������U��p8�P@�Rh]�����������������U��p8�P@�Rl]�����������������U��p8�P@�Rp]�����������������U��p8���   ���   ]�����������U��p8���   ���   ]����������̡p8�P@�Bt����̡p8�P@�Bx�����U��p8�P@�R|]����������������̡p8�P@���   ��p8���   �Bt��U��p8�P@���   ]�������������̡p8�P@���   ��U��p8�P@���   ]��������������U��p8�P@���   ]��������������U��p8�P@���   ]��������������U��p8�P@���   ]��������������U��p8V��H@�QV�ҋM����t��#����p8�Q@P�BV�Ѓ�^]� �̡p8�PH���   Q�Ѓ�������������U��p8�P@�EPQ�JL�у�]� ���̡p8�P@�BHQ�Ѓ����������������U��p8�P@�EP�EP�EPQ�J�у�]� ������������U��p8�P@�EPQ�J�у�]� ����U��p8�P@�EP�EPQ�J�у�]� U��p8�P@�EPQ�J �у�]� ����U��p8���   �R]��������������U��p8���   �R]��������������U��p8���   �R ]��������������U��p8���   ���   ]�����������U��p8���   ��D  ]�����������U��p8�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U��p8���   ���   ]����������̡p8���   �B$��p8�H@�Q0�����U��p8�H@�A4j�URj �Ѓ�]����U��p8�H@�A4j�URh   @�Ѓ�]�U��p8�H@�U�E�I4RPj �у�]�̡p8�H|�������U��V�u���t�p8�Q|P�B�Ѓ��    ^]��������̡p8�H|�Q �����U��V�u���t�p8�Q|P�B(�Ѓ��    ^]��������̡p8�H@�Q0�����U��V�u���t�p8�Q@P�B�Ѓ��    ^]���������U��p8�H@���   ]��������������U��V�u���t�p8�Q@P�B�Ѓ��    ^]��������̡p8�PH���   Q�Ѓ�������������U��p8�PH�EPQ��d  �у�]� �U��p8�H �IH]�����������������U��}qF uHV�u��t?�p8���   �BDW�}W���Ћp8�Q@�B,W�Ћp8�Q�M�Rp��VQ����_^]����������̡p8�P@�BT�����U��p8�P@�RX]�����������������U��p8�P@�R\]����������������̡p8�P@�B`�����U��p8�H��T  ]��������������U��p8�H@�U�A,SVWR�Ћp8�Q@�J,���EP�ыp8�Z��h��hE  �΋��&��Ph��hE  �����P��T  �Ѓ�_^[]����U��p8�PT�EP�EPQ�J�у�]� U��p8�PT�EPQ�J�у�]� ����U��p8�PT�EPQ�J�у�]� ����U��p8�PT�E�R<��PQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��p8�HT�]��U��p8�H@�AV�u�R�Ѓ��    ^]�������������̡p8�HT�hG  �҃�������������U��p8�H@�AV�u�R�Ѓ��    ^]�������������̋�� ����������������������̅�t��j�����̡p8�P��  ��p8�P��(  ��U��p8�P��   ��V�E�P�ҋuP��������M��"�����^��]� ��������̡p8�P��$  ��U��p8�H��  ]��������������U��p8�H���  ]�������������̡p8�H��  ��U��p8�H���  ]��������������U��p8�H��x  ]��������������U��p8�H��|  ]��������������U���EV�����t	V�������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U��p8�H�QV�uV�҃���^]� �3�� �����������3�� �����������U����   h�   ��@���j P�$�  �M�Eh�   ��@���R�M��MPQjǅ`���    ��.���� ��]���U����   V�u��u3�^��]�h�   ��@���j P�Ŋ  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD����l�E�pq�E�`��E����E�0��E� ��E� ��E��q�T.���� ^��]�������������U���   SV�u(3ۉ]���u�p8�H�A�UR�Ѓ�^3�[��]Ëp8�Q�B<W�M3��Ѕ��'  �  �E���tq�MQ�M�����Wh<��M��k���P�M������u�Wj��U�R�E�P��\���Q�_?�E�����P��x���R�U�����P�E�P�H�����P����  �E���t�E� �� t�M�����������t��x������������t��\������������t�M̃��������t�p8�Q�J�E�P����у���t�M��`����}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�  ����E$�M�UVP�Ej QRP����������p8�Q�J�EP�у���_^[��]���������������̋�`����������̋�`����������̡p8�H\�������U��p8�H\�AV�u�R�Ѓ��    ^]�������������̡p8�P\�BQ�Ѓ���������������̡p8�P\�BQ�Ѓ����������������U��p8�P\�EPQ�J�у�]� ����U��p8�P\�EP�EPQ�J�у�]� U��p8�P\�EPQ�J�у�]� ���̡p8�P\�BQ�Ѓ����������������U��p8�P\�EPQ�J �у�]� ����U��p8�P\�EP�EPQ�J$�у�]� U��p8�P\�EP�EP�EPQ�J(�у�]� ������������U��p8�P\�EPQ�J0�у�]� ����U��p8�P\�EPQ�J@�у�]� ����U��p8�P\�EPQ�JD�у�]� ����U��p8�P\�EPQ�JH�у�]� ���̡p8�P\�B4Q�Ѓ����������������U��p8�P\�EP�EPQ�J8�у�]� U��p8�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu������p8�H\�QV�҃���S������3���~=��I �p8�H\�U�R�U��EP�A(VR�ЋM��Q���X����U�R���M���F;�|�_^[��]� ���������������U���VW�}�E��P�������}� ��   �p8�Q\�BV�Ѓ��M�Q���q����E���t]S3ۅ�~H�I �UR���U����E�P���J����E;E�!���p8�Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� �p8�H���   ��U��p8�H���   V�u�R�Ѓ��    ^]����������̡p8�P���   Q�Ѓ�������������U��p8�P�EPQ���   �у�]� ̡p8�H�������U��p8�H�AV�u�R�Ѓ��    ^]��������������U��p8�H�AV�u�R�Ѓ��    ^]��������������U��p8�P��Vh�  Q���   �E�P�ыp8���   �Q8P�ҋ�p8���   ��U�R�Ѓ���^��]��������������̡p8�P�BQ�Ѓ����������������U��p8�P�EPQ�J\�у�]� ����U��p8�P�EP�EP�EP�EP�EPQ���   �у�]� �U��p8�P�EP�EP�EP�EPQ�JX�у�]� �������̡p8�P�B Q��Y�U��p8�P�EP�EP�EP�EPQ���   �у�]� �����U��p8�P�EP�EP�EPQ�J�у�]� ������������U��p8�H��   ]��������������U��p8�P�R$]�����������������U��p8�P��x  ]��������������U��p8�P�EP�EP�EP�EPQ�J(�у�]� ��������U��p8�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U��p8�P�EP�EP�EP�EPQ�J,�у�]� ��������U��p8V��H�QWV�ҋ��p8�H�QV�ҋp8�Q�M�R4Q�MQ�MQOWHPj j V�҃�(_^]� ���������������U��p8�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U��p8�P�EP�EPQ�J@�у�]� U��p8�P�EPQ�JD�у�]� ���̡p8�P�BLQ�Ѓ���������������̡p8�P�BLQ�Ѓ���������������̡p8�P�BPQ�Ѓ����������������U��p8�P�EPQ�JT�у�]� ����U��p8�P�EPQ�JT�у�]� ����U��p8�P�EP�EPQ���   �у�]� �������������U��p8�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �p8���   j P�BV�Ћp8���   �
�E�P�у� ��^��]� ������̡p8�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡p8�H�������U��p8�H�AV�u�R�Ѓ��    ^]��������������U��p8�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U��p8�P�EPQ�J�у�]� ���̡p8�P�BQ��Y�U��p8�P�EP�EPQ�J�у�]� U��VW��������M�U�x@�EPQR��������H ���_^]� �U��VW�������M�U�xD�EPQR�������H ���_^]� �V�������xH u3�^�W���v����΍xH�l����H �_^�����U��V���U����xL u3�^]� W���@����M�U�xL�EPQR���*����H ���_^]� �������������U��V�������xP u���^]� W��������M�U�xP�EP�EQRP��������H ���_^]� ��������U��V�������xT u���^]� W�������M�xT�EPQ�������H ���_^]� U���S�]VW���t.�M��v������_����xL�E�P���Q����H ��ҍM������}��tZ�p8�H�A�U�R�Ћp8�Q�J�E�WP�ыp8�B�P�M�Q�҃���������@@��t�p8�QWP�B�Ѓ�_^[��]� ������U��V��������x` u
� }  ^]� W�������x`�EP�������H ���_^]� ��U��VW�������xH�EP���v����H ���_^]� ���������U��SVW���S����x` u� }  �#���?����x`�E���P���,����H ��ҋ��p8�H�]�QS�҃�;�A�p8�H�QS�҃�;�,��������M�U�xD�EPQSR��������H ���_^[]� _^�����[]� ��������������U��V�������xP u
�����^]� W�������M�U�xP�EP�EQ�MR�UPQR���k����H ���_^]� ��������������U��V���E����xT u
�����^]� W���-����M�xT�EPQ�������H ���_^]� ��������������U��V��������xX tW��������xX�EP��������H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��88  ����t.�E�;�t'�p8�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡p8�H��   ��U��p8�H��$  V�u�R�Ѓ��    ^]�����������U��p8�UV��H��(  VR�Ѓ���^]� �����������U��p8�P�EQ��,  P�у�]� �U��p8�P�EQ��,  P�у����@]� �����������̡p8�H��0  ��p8�H��4  ��p8�H��p  ��p8�H��t  ��U��E��t�@�3��p8�RP��8  Q�Ѓ�]� �����U��p8�P�EPQ��<  �у�]� �U��p8�P�EP�EP�EPQ��@  �у�]� ���������U��p8�P�EP�EPQ��D  �у�]� �������������U��p8�P�EPQ��H  �у�]� �U��p8�P�E��L  ��VWPQ�M�Q�ҋu���p8�H�QV�ҡp8�H�QVW�ҡp8�H�A�U�R�Ѓ�_��^��]� ��������������̡p8�P��T  Q�Ѓ�������������U��p8�P�EPQ��l  �у�]� ̡p8�P��P  Q�Ѓ�������������U��p8�P�EPQ��X  �у�]� ̡p8�H��\  ��U��p8�H��`  V�u�R�Ѓ��    ^]�����������U��p8�P�EP�EP�EP�EP�EPQ��d  �у�]� �U��p8�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���b�����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���o����xP t$S���a���j j �XPj�FP���M����H ���[�    �~` t�p8�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx�p8�Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�T������u#���h���p8�H��0  h�   �҃��E�~P�������j j jW�^����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    �p8�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ������F|��u�E�~x��t�    �F`_^]� �M�Fx������t�3�_^]� U��QVW�}����>[  �p8�H�QhV�҃����p8u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���Y  �EF;u�|�UR�������_�   ^��]� �������������U��QVW�}����~Z  �p8�H�QhV�҃����p8u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'���p8�QP�Bh�Ѓ���t�M��R���,X  F;u�|ʍEP�������_�   ^��]� �������������h��h�   h�8h�   ���������t�������3��������V���(����N^�������������������U��VW�}�7��t��������N�����V�������    _^]�U���EV���V��������Au�p8�H��0  h��j,�����^��^]� �����U���W������G���U�� �������A�  ������A��   �(�������AuR������AuKV���+s  ���$s  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������= ���������Au6�����������U������G�����_��������Au�����U����_�
����������v  �E����U�����������A{���������__��]�������������__��]����U���8�V�E��������At���0�������Au�������������$��p  ���������^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3�����;���W���$���Qp  ��E�����$�<p  �V����������Au�p8�H��0  h��j�����^����_u������������^]� ���U������EV�ы�������z!�p8�؋H��0  h��j5�����U������$�o  �]��F�$�o  �}��$�o  ��E�$�o  �^�����&���^��]� ��������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V������������   �ESP�M�������p8�Q�J�E�P�ыp8�B�Pj j��M�h<�Q�҃��E�P�M�輼��j j��M�Q�U�R��d���P�d�����P�M�Q�w�����P�U�R�j������P��������M��������M�������d����޼���M��ּ���p8�H�A�U�R�Ѓ��M�躼����[t	V��������^��]� ���U��EVP���a��������^]� �����Q�����Y���������U��E�M�U�H4�M�P �U��M�@�l�@8pq�@<�q�@@`��@D ��@H ��@L���@P���@l���@X@��@\��@`@��@d ��@T0��@h0��@p���@t ��P0�H(�@,    ]��������������U���   h�   ��`���j P�Dk  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�����8��]��������������̋�`����������̋�`0����������̋�`@����������̋�`����������̋�`,�����������3�� �����������3�� �����������3�� ���������������������������3�� �����������3��  ����������̸   � ��������3�� �����������3�� ������������ �������������3�� �����������U��P�EQj RPV������M�����   ǆ�   �ǆ�   ��ǆ�   �ǆ�    �ǆ�   @�ǆ�   `�ǆ�    �ǆ�   P�ǆ�   0�ǆ�   P�ǆ�   �]���U���   Vh   ������j P�Ci  �M�U�E Q�MR�U�������7����M�Uh   ��PQRj
�����(^��]��������̋�`\����������̋�`l����������̋�`P����������̋�``����������̋�`T����������̋�`d����������̋�`X����������̋�`h�����������U��p8���   �BXQ�Ѓ���u]� �p8�Q|�M�RQ�MQP�҃�]� ���U��p8���   �BXQ�Ѓ���u]� �p8�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ��p8�Qj j P�B�ЉF����^]� ��̡p8Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� �p8�Q�MP�EP�Q�JP�у��F�   ^]� ����U��E��u�E�M��8��8�   ]� �����������U��EHV����   �$�ȓ�   ^]á�8@��8��uT�EP�'�����=�.  }�����^]Ëu��t�h@�jmh�8j��������t ���-�����8��tV���<����   ^]���8    �   ^]ËM�UQR��|���������H^]�^]�|���-�8u.�|���}�����8��t��謶��V�v�������8    �   ^]Ã��^]ÍI ��y���ؒ��^�U��E�M�UP��P�EjP�����]��������������̸   �����������U��V�u��t���u6�EjP�������u3�^]Ë������t���t��U3�;P��I#�^]�����������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������h�8Ph^� �0������������������U��Vh�8jh^� ���	�������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh�8jh^� �����������t�@��tV�Ѓ�^�3�^���U��Vh�8jh^� ����������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh�8jh^� ���S�������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u���c����N`�[������   �P�����   �E�����ݞ�  ��^��]� ����U��Vh�8jh^� �����������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh�8jh^� ����������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh�8j h^� ���I�������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�8j$h^� �����������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�8j(h^� ����������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh�8j,h^� ���x�������t �@,�E���t�E�MPQV�U���^��]� ��^��]� ��������U��Vh�8j0h^� ���)�������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh�8j4h^� �����������t�@4��tV�Ѓ�^�3�^���Vh�8j8h^� ����������t�@8��tV�Ѓ�^�������U���`Vh�8jDh^� ���v�������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u��������^��]� ����U��Vh�8jHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh�8jLh^� �����������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh�8jPh^� ����������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh�8jTh^� ���Y�������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh�8jXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh�8j`h^� ����������t�@`��tV�Ѓ�^�3�^���U��Vh�8jdh^� ����������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh�8jhh^� ���F�������t1�@h��t*�MQ�U�VR�Ћu��P�������M��������^��]� �u��贆����^��]� �����������Vh�8jph^� �����������t�@p��tV�Ѓ�^Ã��^��Vh�8jlh^� ����������t�@l��tV�Ѓ�^Ã��^��Vh�8jth^� ���|�������t�@t��tV�Ѓ�^�3�^���U��Vh�8jxh^� ���I�������t�@x��t
�MQV�Ѓ�^]� ������������Vh�8j|h^� ����������t�@|��tV�Ѓ�^�������Vh�8h�   h^� �����������t���   ��tV�Ѓ�^�U��Vh�8h�   h^� ����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh�8h�   h^� ���V�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh�8h�   h^� ����������tU���   ��tKW�M�VQ�Ћp8�u���B�HV�ыp8�B�HVW�ыp8�B�P�M�Q�҃�_��^��]� �p8�H�u�QV�҃���^��]� ����������Vh�8h�   h^� ���i�������t���   ��tV�Ѓ�^Ã��^������������U��Vh�8h�   h^� ���&�������t���   ��t
�MQV�Ѓ�^]� ������U��Vh�8h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�8h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh�8h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U��Vh�8h�   h^� ����������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh�8h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh�8h�   h^� ���f�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�8h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�8h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�8h�   h^� ���v�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh�8h�   h^� ���)�������t���   ��tV�Ѓ�^�3�^�������������Vh�8h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������Vh�8h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh�8h�   h^� ���i�������t���   ��tV�Ѓ�^�3�^�������������U��Vh�8h�   h^� ���&�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh�8h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U���Vh�8h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�8h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�8h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U���Vh�8h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�8h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�8h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh�8h�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh�8h�   h^� ���E�������t#���   �E���t�E�MPQV�U���^��]� ��^��]� ��U��Vh�8h�   h^� �����������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh�8h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�8h�   h^� ���V�������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�8h   h^� ����������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh�8h  h^� ����������t��  ��tV�Ѓ�^�3�^�������������U���Vh�8h  h^� ���s�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�8h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�8h  h^� ���s�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh�8h  h^� �����������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�8h  h^� ����������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�8h  h^� ���v�������t��  ��t
�MQV�Ѓ�^]� ������Vh�8h   h^� ���9�������t��   ��tV�Ѓ�^�3�^�������������U��Vh�8h$  h^� �����������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�8h(  h^� ����������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�8h,  h^� ���V�������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�8h0  h^� ���	�������t��0  ��tV�Ѓ�^�3�^�������������U��Vh�8h4  h^� �����������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�8h8  h^� ���v�������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�8h<  h^� ���&�������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh�8h@  h^� �����������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�8hD  h^� ����������t��D  ��tV�Ѓ�^�3�^�������������U��Vh�8hH  h^� ���F�������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�8hL  h^� �����������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�8hP  h^� ����������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh�8hT  h^� ���U�������t'��T  �E���t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh�8hX  h^� �����������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh�8j<h^� ����������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh�8j@h^� ���i�������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h�8Ph�� �0������������������h�8jh�� ��������uË@����U��V�u�> t/h�8jh�� ���������t��U�M�@R�Ѓ��    ^]���U��Vh�8jh�� ����������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�8jh�� ���Y�������t�@��t�M�UQR����^]� ����������U��Vh�8jh�� ����������t�@��t�M�UQR����^]� ����������U��Vh�8jh�� �����������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�8j h�� ����������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�8j$h�� ���9�������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�8j(h�� �����������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�8j,h�� ����������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh�8j0h�� ���9�������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�8j4h�� �����������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh�8j8h�� ����������t�@8�E���t�E�MPQ���U�^��]� ��^��]� ����������U��Vh�8j<h�� ���9�������t�@<��t�M�UQR����^]� ����������U��Vh�8j@h�� �����������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh�8jHh�� ����������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh�8jDh�� ���y�������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh�8jLh�� ���8�������t#�@L�E���t�E�EP�����$�U�^��]� ��^��]� �����U��Vh�8jPh�� �����������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh�8jTh�� ����������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�8jXh�� ���Y�������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�8j\h�� ���	�������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h�8jh�� ��������t�@�ЉF�~��t6h�8jh�� ��������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h�8jh�� �1�������t�@��t�M�UQR���Ѓ~ t1h�8jh�� � �������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h�8jh�� ��������t�@�ЉF�v��t+h�8jh�� ��������t�@��t�M�UQR����^]� �������������U��V�q��t@h�8jh�� �D�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h�8j h�� ���������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h�8jh�� ��������t�@�ЉF�}�]�M�UWSQR���k1  ��t�N��t�E�UWSPR����_^[]� _^3�[]� �U��V�q��t8h�8j(h�� �$�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��I��t)�E$�E�UP�E���\$�E�$R�UPR����]�  3�]�  �������U��V�q��t<h�8j0h�� ��������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��h�8Ph�f �P������������������U��h�8jh�f �,�������t
�@��t]�����]�������U��Vh�8jh�f �����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R躑���E�NP�у�4�M��������^]ÍM�ב�����^]��U��h�8jh�f ��������t
�@��t]��3�]��������U��h�8jh�f �\�������t�x t�P]��3�]������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������A  ����������D�Ez��^�P�P�]��������������N�X�N^�X]���U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��U�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A������������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V�����FP�ޭ��3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  S�]���i  ��؋�U��M�U��U��@�����@�U��@�B�@�������@���@�G�>��w����U���  �w�������F�B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]؋�R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[������E��KH��P�E�SL��H�щKP�P�ST�H�KX�P�����S\��z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����M��}������3�3����u��u�|+�A�����B�4�u�0u��u�p�����u�u�U�E;�}�Q���E����U��U��1���@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���@�D��KX�@�U�����]��C���@�K0���@�KH���C ��C�@�K8���@�KP���C(��C�C@�H���@3����KX���U��r  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������]��E�E����]���E����]��E׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���@�   �KXE)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� ����h�8Ph_� ��������������������h�8jh_� ��������uË@����U��V�u�> t/h�8jh_� �s�������t��U�M�@R�Ѓ��    ^]���U��Vh�8jh_� ���9�������t�@��t�MQ����^]� 3�^]� �������U��Vh�8jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh�8jh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�8jh_� ���i�������t�@��t�MQ����^]� 3�^]� �������U��Vh�8j h_� ���)�������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�8j$h_� �����������t�@$��t�MQ����^]� 2�^]� �������Vh�8j(h_� ����������t�@(��t��^��3�^������Vh�8j,h_� ���|�������t�@,��t��^��3�^������U��Vh�8j0h_� ���I�������t�@0��t�MQ����^]� 3�^]� �������U��Vh�8j4h_� ���	�������t�@4��t�M�UQR����^]� ���^]� ��Vh�8j8h_� �����������t�@8��t��^��3�^������U��Vh�8j<h_� ����������t�@<��t�MQ����^]� ��������������U��Vh�8j@h_� ���Y�������t�@@��t�MQ����^]� ��������������U��Vh�8jDh_� ����������t�@D��t�MQ����^]� 3�^]� �������U��Vh�8jHh_� �����������t�@H��t�MQ����^]� ��������������Vh�8jLh_� ����������t�@L��t��^��3�^������Vh�8jPh_� ���l�������t�@P��t��^��3�^������Vh�8jTh_� ���<�������t�@T��t��^��^��������Vh�8jXh_� ����������t�@X��t��^��^��������Vh�8j\h_� �����������t�@\��t��^��^��������U��Vh�8j`h_� ����������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�8jdh_� ���i�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh�8jhh_� ���)�������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�8jlh_� �����������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�8jph_� ����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�8jth_� ���I�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�8jxh_� ���	�������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh�8j|h_� �����������t�@|��t�MQ����^]� 3�^]� �������U��Vh�8h�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�8h�   h_� ���6�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�8h�   h_� ���ֿ������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�8h�   h_� ���v�������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U��������������������x*  ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@����A���E�    �����]����]��]�����������]����]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�����F�@��R�M������~���Q�M��y����v;�t�v��P�M��c����M����m��M�u�_^[�M�UQR�M�������]� ����������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$����E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��2�H�[�o�������U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V藖���FP莖��3����F�F^��U��SV��WV�r����^S�i����E3����~�~;�t_�p8�Q���   h����jIP�у��;�t9�}��t;�p8�B���   h����    jNQ�҃����uV�������_^3�[]� �E�~_�F^�   []� ����������U��SV��WV����^S蹕���}3Ƀ��N�N;���   9��   �G;���   �p8�Q���  h����jlP�у����t=� t@�G��t9�p8�Jh����    ���  jqR�Ѓ����u���=���_^3�[]� �O�N�G�Q��    R�F�QP�  �����t�N�WP��QPR�x  ��_^�   []� ���������U��SV��WV����~W蹔��3Ƀ��N�N9M��   �E;���   ��    �p8�H���  h��h�   S�҃����t=�} tH�E��tA�p8�Q���  h����h�   P�у����u���B���_^3�[]� �U�V�,�F   �p8�H���  h��h�   j�҃����t��E�M�F�PSPQ�q  �E����t!�V�?�W�RWP�U  ��_^�   []� ��M�_^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��S�]V��3�W�~���F�F�CV;C��   ����W�����3��F�F�p8�Q���   h��jIj�Ѓ������   �p8�Q���   h��jNj�Ѓ����uV覒����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �`���W�Z���3��F�F�p8�B���   h��jIj�у����t[�p8�B���   h��jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�`  ��]������������V��FW��u�~��N�<��u�< ��u_3�^áp8�H�F��  h��j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�#���3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�(��-���3����_�F�F^��������������U���SV�uW���^S�}������3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY�p8�H���  h��j8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E�0��k�����]� �����U����Q�Ej�E��A�MRPQ�M��E�0�������]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�����t!�A��t�B�A�Q�P�A    �A    �̋�� 8��@���HV3��q�q�P�r�r����p�p�p�P�H^������V���8������F3��F��;�t�N;�t�H�F�N�H�V�V�F�F��;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3����;�t�F;�t�A�F�N�H�V�V�Et	V��������^]� ������������U��V��W�~W�(��z���3����E��F�Ft	V行����_��^]� ������U��V��������Et	V�y�������^]� ���������������U��p8�PH�EPQ���  �у�]� �U��p8�P�B4VW�}j��h�  ���ЋMWQ���D  _^]� ��������������U��V���PXW�ҋ}P���'=�����Et�_�   ^]� �M�UPWQR���1  _^]� �����������U��S�]VW��j ����:���8�  �}uI�~ uC�p8�P���   j h�  ���Ѕ�u�p8�QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ����  _^[]� ��������U��EP�A    ������]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �}  ����   �M3�V�
:���8�  u4����P�w蔮���p8�P�M�B4��jh�  ��_^�C�[��]� �MV��9���8�  u�E�M��RPQ����_^�   [��]� �MV�9���8�  t�MV�9���8��  �p8�P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P����3��؃��u�;�t�p8�QH���  VS�Ѓ��E��M�;O�f  9w�]  �p8�B�M���   Vh�  �҅�u!�p8�P�M���   Vh�  �Ѕ��  �p8�Q�M�B4Vh�  ��;�t
V���������E��G�p8���   ���   �Ћ]�E�;���   ;���   S�7����M���jQ�ˉu��uĉuȉủuЉu؉u������U�E��ˉu��u�u�U�E��]��E�   ������t!��t��t�u���E�   ��E�   ��E�   �:����M�;�t�N�����BX�M�Q����P�����M܃�;�t�L����M��T����M��L����M������]�M�U�EQSRP����  _^[��]� �M�����_^�   [��]� �������������̸   � ��������� ������������̃��� ����������� �������������U��p8�H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� �p8�Q0�F�M���   PQW�ҋF��^_]� U��p8�H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U��p8�H���  ]��������������U��p8�H���  ]��������������U��p8�P�EP�EP�EP�EPQ���   �у�]� �����U��p8�E�P�EP�E���\$�E�$PQ���   �у�]� �������������U��p8�P�EP�EP�EPQ���   �у�]� ��������̡p8�P���   Q�Ѓ�������������U��p8�P�EP�EP�EPQ���   �у�]� ���������U��p8�P�EP�EPQ���   �у�]� �������������U��p8�H�U�ApR�Ѓ�]� �����U��p8�P�EP�EPQ���  �у�]� �������������U��p8�P�EP�EPQ���  �у�]� �������������U��p8�P�EP�EPQ���  �у�]� �������������U��p8�P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P�	  ��R���E�P���ҡp8�P�B<�M��Ћ}��t0j �M�QW��G������u�p8�B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4����l�E����E����E�0��E�@��E���E�pq�E��qǅx���`�ǅ|��� ��E� ��E�@��E����E���E�P��E����E���E�0��E� ��E����E�0��X����p8���B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u�p8�H�A�UR�Ѓ�^3�[��]Ëp8�Q�B<W�M3��Ѕ��'  范���E���tq�MQ�M��W��Wh<��M��[��P�M��W���u�Wj��U�R�E�P��\���Q�_?�5k����P��x���R�E[����P�E�P�8[����P���̈́���E���t�E� �� t�M�����W����t��x�������W����t��\�������W����t�M̃���zW����t�p8�Q�J�E�P����у���t�M��PW���}� t"�U(�E$�M�R�UP�EQ�MRPQ���������U�R��������E$�M�UVP�Ej QRP����������p8�Q�J�EP�у���_^[��]����������������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`<����������̋�`L����������̋�` ����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`����������̋�`(����������̋�`8����������̋�`H����������̋�`����#��#���#4��#m��#���#��#��#���#T��#�Ë�U�������r  �} ��8t��  ��]Ë�Q�L��y  YË�U��V��������EtV���Y��^]� ��U��EVW��u|P�*  Y��u3��  �  ��u�*  ���"*  ����T��(  ��8��"  ��}�   ���(  ��| �%  ��|j �   Y��u��8�   �%  ��3�;�u19=�8~���89=9u�C"  9}u{��$  �  �*  �j��uY�y  h  j��  ��YY;��6���V�5�#�5�8��  Y�Ѕ�tWV�  YY� ��N���V�7  Y�������uW�4  Y3�@_^]� jh��+  ����]3�@�E��u9�8��   �e� ;�t��u.�P���tWVS�ЉE�}� ��   WVS�r����E����   WVS�֛���E��u$��u WPS���Wj S�B����P���tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�P���tWVS�ЉE��E������E���E��	PQ�*  YYËe��E�����3���*  Ë�U��}u�x,  �u�M�U�����Y]� ��U��QSVW�5�T�h  �5�T���}��X  ��YY;���   ��+ߍC��rwW�,  ���CY;�sH�   ;�s���;�rP�u��7  YY��u�G;�r@P�u��!  YY��t1��P�4��s  Y��T�u�e  ���V�Z  Y��T�EY�3�_^[�Ë�Vjj �  ��V�3  ����T��T��ujX^Ã& 3�^�jh��)  �  �e� �u�����Y�E��E������	   �E��)  ��j  Ë�U���u���������YH]��5L=�3  Y��t��j�-  jj �U-  ���6,  jh��	)  �e� �u;5�Sw"j�0  Y�e� V��8  Y�E��E������	   �E��)  �j�/  YË�U��V�u�����   SW�=��=,: u�.  j��,  h�   �  YY��S��u��t���3�@P���uV�S���Y��u��uF�����Vj �5,:�׋؅�u.j^9�>t�u�;  Y��t�u�{����#;  �0�;  �0_��[�V�f;  Y�;  �    3�^]��������̋T$�L$��ti3��D$��u��   r�=�S t�;  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh �n'  �u��tu�=�SuCj�/  Y�e� V�G/  Y�E��t	VP�h/  YY�E������   �}� u7�u�
j�.  Y�Vj �5,:����u�:  ����P�9  �Y�2'  �;@#u����<  ��������̃=�S ��@  ���\$�D$%�  =�  u�<$f�$f��f���d$�V@  � �~D$f(p�f(�f(�fs�4f~�fT��f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�=  ���D$��~D$f��f(�f��=�  |!=2  �fT`��\�f�L$�D$����f���fV��fT��f�\$�D$���������������̃=�S t-U�������$�,$�Ã=�S t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�������U��WV�u�M�}�����;�v;���  ��   r�=�S tWV����;�^_u^_]��?  ��   u������r*��$�d���Ǻ   ��r����$�x��$�t���$����������#ъ��F�G�F���G������r���$�d��I #ъ��F���G������r���$�d��#ъ���������r���$�d��I [�H�@�8�0�(� ���D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�d���t�|������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�  �����$����I �Ǻ   ��r��+��$���$�  ��8�`��F#шG��������r�����$�  �I �F#шG�F���G������r�����$�  ��F#шG�F�G�F���G�������V�������$�  �I �����������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�  ��  ( < �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̺P#�>  �P#�|=  �Ƀ=�8t�����K  �����z�����������������̃��$�P  �   ��ÍT$�O  R��<$�D$tQf�<$t�pO  �   �u���=�8 ��O  �   ��#��O  �  �u,��� u%�|$ u���EO  �"��� u�|$ u�%   �t����-�'�   �=�8 ��O  �   ��#�N  ZË�U��EV���F ��uc�  �F�Hl��Hh�N�;8/t�T.�Hpu��Y  ��F;X-t�F�T.�Hpu�YR  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P��\  ��e�F�P�[  ��Yu��P��\  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�\  �M��E��M��H��EP�\  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�`  @PV�V�]  ��^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+�/1  j_VVVVV�8�gY  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	��0  j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h��SV��_  ��3ۅ�tSSSSS�xW  ���N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�Bt�90uj�APQ�[  ���}� t�E��`p�3�_^[�Ë�U���,�@#3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�a  3ۃ�;�u�/  SSSSS�0��W  �����o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�4_  ��;�t���u�E�SP�u��V�u��������M�_^3�[�(����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �C���9}}�}�u;�u+�.  j^WWWWW�0��V  ���}� t�E�`p����  9}vЋE��� 9Ew	�|.  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV��J  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� ��_  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �_  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�q�����u�E�8 u���} �4����$�p���WF�_  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��]  0�F�U�����;�u��|��drj jdRP��]  0��U�F����;�u��|��
rj j
RP�]  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�������u-�Y+  j^�03�PPPPP�S  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�������}� t�E��`p�3�_^[�Ë�U���,�@#3ŉE��ESVW�}j^V�M�Q�M�Q�p�0��[  3ۃ�;�u�J*  SSSSS�0�R  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P��Y  ��;�t���u�E�SV�u���`������M�_^3�[������Ë�U���0�@#3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�[  3ۃ�;�u�)  SSSSS�8��Q  �����   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW�4Y  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[������Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����#�6�  ��Y���(r�_^Ë�Vh   h   3�V��Z  ����tVVVVV�O  ��^Ë�U�������]�����]��E��u��M��m��]����]�����z3�@��3���h������th��P����tj �������jh �i  j�*  Y�e� �u�N��t/��8��8�E��t9u,�H�JP����Y�v����Y�f �E������
   �X  Ë���j��  Y�̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U��V�5�#�5 ��օ�t!��#���tP�5�#���Ѕ�t���  �'� �V����uV�  Y��th��P����t�u�ЉE�E^]�j ����YË�U��V�5�#�5 ��օ�t!��#���tP�5�#���Ѕ�t���  �'� �V����uV�   Y��th�P����t�u�ЉE�E^]��$�� ��V�5�#� �����u�5�8�e���Y��V�5�#�(���^á�#���tP�5�8�;���Y�Ѓ�#���#���tP�,���#��  jh@�	  � �V����uV�a  Y�E�u�F\��3�G�~��t$h��P���Ӊ��  h��u��Ӊ��  �~pƆ�   CƆK  C�Fh0)j�`  Y�e� �vh�0��E������>   j�?  Y�}��E�Fl��u�8/�Fl�vl�I  Y�E������   �  �3�G�uj�'  Y�j�  YË�VW���5�#�������Ћ���uNh  j��  ��YY��t:V�5�#�5�8�����Y�Ѕ�tj V�����YY� ��N���	V�J���Y3�W�4�_��^Ë�V��������uj�>  Y��^�jhh�  �u����   �F$��tP�����Y�F,��tP�����Y�F4��tP�����Y�F<��tP�����Y�F@��tP�����Y�FD��tP����Y�FH��tP����Y�F\=��tP����Yj��  Y�e� �~h��tW�8���u��0)tW�k���Y�E������W   j�  Y�E�   �~l��t#W�H  Y;=8/t��`.t�? uW�F  Y�E������   V����Y��  � �uj�h  YËuj�\  YË�U��=�#�tK�} u'V�5�#�5 ��օ�t�5�#�5�#���ЉE^j �5�#�5�8����Y���u�x�����#���t	j P�(�]Ë�VW� �V����uV�R  Y�����^  �5�hL�W��h@�W��8��h4�W��8��h,�W��8�փ=�8 �5(���8t�=�8 t�=�8 t��u$� ���8�,���8U�5�8��8�$���#�����   �5�8P�օ���   �_  �5�8�����5�8��8�����5�8��8�����5�8��8�u�������8�0  ��tehI�5�8�����Y�У�#���tHh  j�   ��YY��t4V�5�#�5�8����Y�Ѕ�tj V�y���YY� ��N��3�@��$���3�_^Ë�U��VW3��u������Y��u'9�8vV�<����  ;�8v��������uʋ�_^]Ë�U��VW3�j �u�u��T  ������u'9�8vV�<����  ;�8v��������uË�_^]Ë�U��VW3��u�u�U  ��YY��u,9Et'9�8vV�<����  ;�8v��������u���_^]Ë�U��W��  W�<��u�����  ��`�  w��t�_]Ë�U���\  �u�  �5�#�D���h�   �Ѓ�]Ë�U��hh�����thX�P����t�u��]Ë�U���u�����Y�u�@��j�  Y�j��  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=<� th<��W  Y��t
�u�<�Y�O���h@�h(�����YY��uBh��������$$��c����=�T Yth�T�V  Y��tj jj ��T3�]�jh��  j��  Y�e� 3�C99��   �9�E�9�} ��   �5�T�����Y���}؅�tx�5�T����Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5�T�~������5�T�q�����9}�u9E�t�}�}؉E����u܋}��hP��D��_���YhX��T��O���Y�E������   �} u(�9j�  Y�u�����3�C�} tj��  Y��8
  Ë�U��j j�u�������]�jj j ������Ë�V������V�  V�kX  V��C  V��  V�JX  V�2V  V�  V�V  h�������$��#^�jTh��s	  3��}��E�P�P��E�����j@j ^V�&���YY;��  ��S�5�S��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@��S��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M����S���S ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=�S|���=�S�e� ��~m�E����tV���tQ��tK�uQ�L���t<�u���������4��S�E� ���Fh�  �FP��V  YY����   �F�E�C�E�9}�|�3ۋ���5�S����t���t�N��r�F���uj�X�
��H������P�H������tC��t?W�L���t4�>%�   ��u�N@�	��u�Nh�  �FP�4V  YY��t7�F�
�N@�����C���g����5�S�D�3��3�@Ëe��E���������q  Ë�VW��S�>��t1��   �� t
�GP�T����@   ;�r��6�u����& Y�����T|�_^Ã=�T u�=  V�5�8W3���u����   <=tGV�H  Y�t���u�jGW�n�����YY�=�8��tˋ5�8S�BV�yH  ��C�>=Yt1jS�@���YY���tNVSP��H  ����t3�PPPPP�i@  �����> u��5�8�����%�8 �' ��T   3�Y[_^��5�8�����%�8 ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�U  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�6T  Y��t��M�E�F��M��E���T  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9�Tu�;  h  � 9VS�$:�X���T�59;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�q�����Y;�t)�U��E�P�WV�}�������E���H��8�5�83�����_^[�Ë�U��(:��SV�5l�W3�3�;�u.�֋�;�t�(:   �#����xu
jX�(:��(:����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5h�SSS+�S��@PWSS�E��։E�;�t/P����Y�E�;�t!SS�u�P�u�WSS�օ�u�u��l���Y�]��]�W�d����\��t;�u��`���;��r���8t
@8u�@8u�+�@P�E��0�����Y;�uV�\��E����u�VW������V�\���_^[�Ë�V����W��;�s���t�Ѓ�;�r�_^Ë�V����W��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P�p��,:��u]�3�@��S]Ã=�SuWS3�9�SW�=�~3V�5�S��h �  j �v��x��6j �5,:�׃�C;�S|�^�5�Sj �5,:��_[�5,:�t��%,: �Ë�U��QQV�G��������F  �V\�@$W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   �4$�=8$���;�}$k��~\�d9 �=4$�8$B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]���h@"d�5    �D$�l$�l$+�SVW�@#1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���̋�U���S�]V�s35@#W��E� �E�   �{���t�N�38�����N�F�38�o����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���xF  �E���|@G�E��؃��u΀}� t$����t�N�38������N�V�3:������E�_^[��]��E�    �ɋM�9csm�u)�=�S t h�S�3J  ����t�UjR��S���M�F  �E9Xth@#W�Ӌ��F  �E�M��H����t�N�38�i����N�V�3:�Y����E��H���E  �����9S�R���h@#W����E  ������U����@#�e� �e� SW�N�@��  ��;�t��t	�УD#�`V�E�P����u�3u����3�� �3����3��E�P�|��E�3E�3�;�u�O�@����u������5@#�։5D#^_[��jh��v���3��]3�;���;�u�b  �    WWWWW�8  ������S�=�Su8j�  Y�}�S�*  Y�E�;�t�s���	�u���u��E������%   9}�uSW�5,:��������6����3��]�u�j��  YË�U���(  �@#3ŉE��D$Vtj
�  Y�I  ��tj�I  Y�D$��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P��������������(�����0���j ǅ����  @��������,��������(���P���j�����̋�U��M�D$�U#U��#�ʉD$]Ë�U��QQS�]VW3�3��}�;�H$t	G�}���r���w  j�M  Y���4  j�M  Y��u�=�8�  ���   �A  h���  S�0:W�=  ����tVVVVV�;5  ��h  �I:Vj �M; �X���u&h��h�  V�q=  ����t3�PPPPP��4  ��V��<  @Y��<v8V�<  ��;�j�D=h��+�QP�L  ����t3�VVVVV�4  ���3�h��SW�xK  ����tVVVVV�4  ���E��4�L$SW�SK  ����tVVVVV�k4  ��h  hX�W��I  ���2j��H���;�t$���tj �E�P�4�L$�6�<  YP�6S���_^[��j�L  Y��tj�L  Y��u�=�8uh�   �)���h�   ����YYË�U��E�L=]Ë�VW3��P=�<�%u�� %�8h�  �0���JH  YY��tF��$|�3�@_^Ã$� % 3����S�T�V� %W�>��t�~tW��W������& Y���� &|ܾ %_���t	�~uP�Ӄ��� &|�^[Ë�U��E�4� %���]�jh������3�G�}�3�9,:u�����j�,���h�   ����YY�u�4� %9t���nj�=���Y��;�u�  �    3��Qj
�Y   Y�]�9u,h�  W�AG  YY��uW�����Y�m  �    �]���>�W�����Y�E������	   �E������j
�(���YË�U��EV�4� %�> uP�"���Y��uj����Y�6���^]Ë�U���S��Sk����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ��>����   ��S�5x�h @  ��H� �  SQ�֋�S��>�   ���	P��>�@��S����    ��>�@�HC��>�H�yC u	�`���>�x�ueSj �p�֡�>�pj �5,:����S��>k���S+ȍL�Q�HQP�3  �E����S;�>v�m��S��S�E��>�=�S[_^�á�SV�5�SW3�;�u4��k�P�5�SW�5,:���;�u3��x��S�5�S��Sk�5�Sh�A  j�5,:���F;�t�jh    h   W����F;�u�vW�5,:��뛃N��>�~��S�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U�����S�Mk��S������M���SI�� VW}�����M���������3���U���S����S�;#U�#��u
���];�r�;�u��S��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1��S�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t��S�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;�>u�M�;�Su�%�> �M���B_^[�Ë�U��E3�;� &tA��-r�H��wjX]Ë�$&]�D���jY;��#���]��������u��'Ã��������u��'Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E��>]Ë�U���5�>����Y��t�u��Y��t3�@]�3�]�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh�����e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E�����Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[��������S3�Ë�U��� S3�9]u �����SSSSS�    ��%  ������   �MV�u;�t!;�u����SSSSS�    ��%  ������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u���>  ����;�t�M�x�E����E�PS�<  YY��_^[�Ë�U���uj �u�u�u�5�����]Ë�U���(  ��?��?��?��?�5�?�=�?f��?f��?f��?f��?f�%�?f�-�?���?�E ��?�E��?�E��?�������?  ��?��>��>	 ���>   �@#�������D#���������� ?j�jI  Yj ���h������= ? uj�FI  Yh	 ����P����Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9�At�5�S�����Y����M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E܄���M��]�Q��]���]���Y����  �1���� "   �  �E܀���M��]�Q��E�   �]���]���Y�j  �E�   �E܀���E�x���]���]���"  �M��E�x��r����E�t��׉M��E�t��Z����E܄�놃�tNIt?It0It ��t����   �E�l���E�d���E܄�����E܄��x����E�   ��������   �E�   �E�\���������������   �$�\;�E�t���E�x���E܀���E�T���E�L���E�D��y����E�<��m����E�8���E�4���E�0���M����]���]�M��]�Q�E�   ��Y��u����� !   �E��_^[���:�:�:�:�:�:{:�:e:\:;;;�%�S �������S3�Ë�U��QQSV���  V�5�'��N  �EYY�M�ظ�  #�QQ�$f;�uU�~M  YY��~-��~��u#�ESQQ�$j� L  ���rVS�N  �EYY�d�ES������\$�E�$jj�?��L  �]��EY�]�Y����DzVS�JN  �E�YY�"�� u��E�S���\$�E�$jj��K  ��^[��U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]��������������U���0���S�ٽ\�����=X/ t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=X/ t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=�8 uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��������������������s4����,ǅr���   ��������������������v���VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�K  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^�����'�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����'�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����'���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�'��p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t��������' u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t��'����'���l$�����'����'���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ��������'�|$�l$�ɛ�l$������l$��Ã�,��?�$�.(����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������' �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����(�Ƀ�u�\$0�|$(���l$�-$(�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�(�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���(�|$�(�<$� �|$$�D$$   �D$(�l$(���(�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������' �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����(�Ƀ�u�\$0�|$(���l$�-$(�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�(�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���(�|$�(�<$� �|$$�D$$   �D$(�l$(���(�<$�l$$�Q�����0Z�����0Z�������@���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�y;  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z����������������������   s��������������������������   v���������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP轧��3��ȋ��~�~�~����~����0)���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �@#3ŉE�SW������P�v����   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�������C�C��u�j �v�������vPW������Pjj �K?  3�S�v������WPW������PW�vS�,=  ��DS�v������WPW������Ph   �vS�=  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[������jh0������������T.�Gpt�l t�wh��uj �>���Y��������j�X���Y�e� �wh�u�;5X-t6��tV�8���u��0)tV����Y�X-�Gh�5X-�u�V�0��E������   뎋u�j����YË�U���S3�S�M�菬����A���u��A   ���8]�tE�M��ap��<���u��A   ����ۃ��u�E��@��A   ��8]�t�E��`p���[�Ë�U��� �@#3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�`-��   �E��0=�   r����  �p  ����  �d  ��P������R  �E�PW������3  h  �CVP����3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�ӣ���M��k�0�u���p-�u��*�F��t(�>����E���\-D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C��d-Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95�A�X�������M�_^3�[������jhP������M���������}�������_h�u�u����E;C�W  h   ����Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�8���u�Fh=0)tP�¢��Y�^hS�=0����Fp��   �T.��   j�����Y�e� �C��A�C��A�C��A3��E��}f�LCf�E�A@��3��E�=  }�L��P+@��3��E�=   }��  ��X,@���5X-�8���u�X-=0)tP�	���Y�X-S���E������   �0j�R���Y��%���u ��0)tS�ӡ��Y�H����    ��e� �E��x���Ã=�T uj��V���Y��T   3�Ë�U��SV�u���   3�W;�to=X1th���   ;�t^9uZ���   ;�t9uP�Z������   �m;  YY���   ;�t9uP�9������   �;  YY���   �!������   ����YY���   ;�tD9u@���   -�   P��������   ��   +�P�������   +�P�Ԡ�����   �ɠ�������   �=�0t9��   uP��8  �7袠��YY�~P�E   ��X.t�;�t9uP�}���Y9_�t�G;�t9uP�f���Y���Mu�V�W���Y_^[]Ë�U��SV�50�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�X.t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�58�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�X.t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu��`.tV�Y���Y��^�3��jhp�Y���蟵����T.�Fpt"�~l t舵���pl��uj �͹��Y���l����j�����Y�e� �Fl�=8/�i����E��E������   ��j�����Y�u�Ë�U��E�B]Ë�U���(  �@#3ŉE������� SjL������j P违����������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   ���������j �������(���P�����u��uj�%  Yh ����P����M�3�[�Ν���Ë�U���5B觱��Y��t]��j��$  Y]������U����u�M�������E����   ~�E�Pj�u�18  ������   �M�H���}� t�M��ap��Ë�U��=�A u�E�(/�A��]�j �u����YY]Ë�U���SV�u�M��t����]�   ;�sT�M胹�   ~�E�PjS�7  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P��7  YY��t�Ej�E��]��E� Y��]���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�1  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=�A u�E�H���w�� ]�j �u�����YY]Ë�U���(�@#3ŉE�SV�uW�u�}�M��"����E�P3�SSSSW�E�P�E�P��A  �E�E�VP�V7  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�@����Ë�U���(�@#3ŉE�SV�uW�u�}�M��z����E�P3�SSSSW�E�P�E�P�CA  �E�E�VP��;  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[蘚������������������U��WV�u�M�}�����;�v;���  ��   r�=�S tWV����;�^_u^_]�I�����   u������r*��$��a��Ǻ   ��r����$��`�$��a��$�xa�a4aXa#ъ��F�G�F���G������r���$��a�I #ъ��F���G������r���$��a�#ъ���������r���$��a�I �a�a�a�a�a�a�a�a�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��a���a�abb�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��c�����$�0c�I �Ǻ   ��r��+��$��b�$��c��b�b�b�F#шG��������r�����$��c�I �F#шG�F���G������r�����$��c��F#шG�F�G�F���G�������V�������$��c�I 4c<cDcLcTc\cdcwc�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��c���c�c�c�c�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��MS3�VW;�t�};�w�]���j^�0SSSSS���������0�u;�u��ڋъ�BF:�tOu�;�u��"���j"Y�����3�_^[]Ë�U��MSV�u3�W�y;�u�����j^�0SSSSS�.��������   9]v݋U;ӈ~���3�@9Ew����j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�a���@PWV�������3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0�@#3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��A  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�<������M�_�s^��3�[�������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j蜭��YË�U��E�M%����#�V������t1W�}3�;�tVV�qJ  YY������j_VVVVV�8� �������_��uP�u��t	�AJ  ���8J  YY3�^]�SVW�T$�D$�L$URPQQh�hd�5    �@#3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C��N  �   �C��N  �d�    ��_^[ËL$�A   �   t3�D$�H3������U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�7N  3�3�3�3�3���U��SVWj j h�iQ�m  _^[]�U�l$RQ�t$������]� jh��1����M3�;�v.j�X3���;E�@u�����    WWWWW�L�����3���   �M��u;�u3�F3ۉ]���wi�=�SuK������u�E;�Sw7j脿��Y�}��u����Y�E��E������_   �]�;�t�uWS蛏����;�uaVj�5,:����;�uL9=�>t3V����Y���r����E;��P����    �E���3��uj�(���Y�;�u�E;�t�    ���e����jh������]��u�u�>���Y��  �u��uS�w���Y�  �=�S��  3��}�����  j葾��Y�}�S躾��Y�E�;���   ;5�SwIVSP��������t�]��5V�k���Y�E�;�t'�C�H;�r��PS�u�聑��S�j����E�SP萾����9}�uH;�u3�F�u������uVW�5,:���E�;�t �C�H;�r��PS�u��-���S�u��C������E������.   �}� u1��uF������uVSj �5,:�������u�]j�¼��YË}����   9=�>t,V����Y�����������9}�ul����P�W���Y��_����   ����9}�th�    �q��uFVSj �5,:�������uV9�>t4V����Y��t���v�V����Y�;����    3��r�����(����|�����u��������P������Y���ҋ�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�h@"d�    P��SVW�@#1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh�諳�������@x��t�e� ���3�@Ëe��E�����襶���ĳ���h-n�����Y�\BË�U��E�`B�dB�hB�lB]Ë�U��E�@$V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5hB����Y�j h�����3��}�}؋]��Lt��jY+�t"+�t+�td+�uD襡�����}؅�u����a  �`B�`B�`�w\���]���������Z�Ã�t<��t+Ht�����    3�PPPPP�������뮾hB�hB��dB�dB�
�lB�lB�E�   P�H����E�Y3��}���   9E�uj�;���9E�tP����Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.�4$�M܋8$�4$�9M�}�M�k��W\�D�E���谞����E������   ��u�wdS�U�Y��]�}؃}� tj �x���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�衱��Ë�U��E�tB]Ë�U��E�xB]�jh0�1����e� �u�u����E��/�E� � �E�3�=  �����Ëe�}�  �uj�4��e� �E������E��#���Ë�U����u�M��@����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U���SVW�X����e� �=|B ����   h� ��������*  �5�h� W�օ��  P袜���$� W�|B��P荜���$� W��B��P�x����$� W��B��P�c���Y��B��th� W��P�K���Y��B��B;�tO9�BtGP詜���5�B��蜜��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9��B;�t0P�Y���Y��t%�ЉE���t��B;�tP�<���Y��t�u��ЉE��5|B�$���Y��t�u�u�u�u����3�_^[�Ë�U��ES3�VW;�t�};�w�����j^�0SSSSS�%��������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u�����j"Y����3�_^[]Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�d���j^�0SSSSS����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x���������j"Y���낋�U��MV3�;�|��~��u��8�(��8��8�����VVVVV�    ����������^]Ë�U��E��t���8��  uP�����Y]Ë�U��QV�uV�O  �E�FY��u�V���� 	   �N ����/  �@t�;���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�iM  �� ;�t�]M  ��@;�u�u��L  Y��uV�L  Y�F  W��   �F�>�H��N+�I;��N~WP�u�K  ���E��M�� �F����y�M���t���t������������S���#�@ tjSSQ��B  #����t%�F�M��3�GW�EP�u�K  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u脾���8*u�ϰ?�d����} �^[]Ë�U���x  �@#3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������z�����u5������    3�PPPPP�1����������� t
�������`p������
  �F@u^V��L  Y��#���t���t�ȃ���������S����A$u����t���t�ȃ�������S����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw���� ��3��3�3���� j��Y������;���	  �$����������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������V  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u�T/������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�J  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  �P/������P����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������G  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�#���������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5�#����Y�Ћ���������   t 9�����u������PS�5�#����Y��YY������gu;�u������PS�5�#�Ȑ��Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�6  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u�P/�������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�D  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t��������x�������� Y���������������t������������������������� t
�������`p��������M�_^3�[�
y���Ð�y�w-x�x�x�x(yVz�%�S �3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u����M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M����X0��{L�H��M�����{,�X0�2��M�����z�X0���M�����z�H0��H0��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E������S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�Э��� "   ]��í��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���`/;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�U�������uV�,���Y�E�^�Ë�d/�h��  �u(�  �u�����E ���Ë�U��=X/ u(�u�E���\$���\$�E�$�uj�/�����$]�謬��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   �@#3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=X/ u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3���q����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-p0�]���t����-p0�]�������t
�-|0�]����t	�������؛�� t���]����jhP�����3�9�StV�E@tH9�0t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�0 �e��U�E�������e��U衖��Ë�S��QQ�����U�k�l$���   �@#3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|������������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�y�����h��  ��x��������>YYt�=X/ uV�q���Y��u�6�I���Y�M�_3�^�7n����]��[Ë�U����@#3ŉE�SV3�W��9�Bu8SS3�GWh�h   S�����t�=�B�����xu
��B   9]~"�M�EI8t@;�u�����E+�H;E}@�E��B����  ;���  ����  �]�9] u��@�E �5��3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�*  ��;�t� ��  �P�Hk��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5��SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�O)  ��;�tj���  ���P�j��Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�����t"SS9]uSS��u�u�u�VS�u �h��E�V�_���Y�u��V����E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�6  Y�E���u3��!  ;E ��   SS�MQ�uP�u ��6  ���E�;�tԋ5��SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�9(  ��;�t����  ���P�pi��Y;�t	� ��  �����3�;�t��u�SW� j�����u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��6  ���u������#u�W�4���Y��u�u�u�u�u�u�����9]�t	�u��%j��Y�E�;�t9EtP�j��Y�ƍe�_^[�M�3��j���Ë�U����u�M���p���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ�@#3ŉE���BSV3�W��;�u:�E�P3�FVh�V�����t�5�B�4����xu
jX��B���B����   ;���   ����   �]�9]u��@�E�5��3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�R&  ��;�t� ��  �P�g��Y;�t	� ��  ���؅�ti�?Pj S�>h����WS�u�uj�u�օ�t�uPS�u����E�S�p����E�Y�u3�9]u��@�E9]u��@�E�u��3  Y���u3��G;EtSS�MQ�uP�u��3  ����;�t܉u�u�u�u�u�u�����;�tV�h��Y�Ǎe�_^[�M�3��h���Ë�U����u�M���n���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v�g���v�g���v�g���v�g���v�g���v�{g���6�tg���v �lg���v$�dg���v(�\g���v,�Tg���v0�Lg���v4�Dg���v�<g���v8�4g���v<�,g����@�v@�!g���vD�g���vH�g���vL�	g���vP�g���vT��f���vX��f���v\��f���v`��f���vd��f���vh��f���vl��f���vp��f���vt�f���vx�f���v|�f����@���   �f�����   �f�����   �f�����   �zf�����   �of�����   �df�����   �Yf�����   �Nf�����   �Cf�����   �8f�����   �-f����,^]Ë�U��V�u��t5�;X1tP�
f��Y�F;\1tP��e��Y�v;5`1tV��e��Y^]Ë�U��V�u��t~�F;d1tP��e��Y�F;h1tP�e��Y�F;l1tP�e��Y�F;p1tP�e��Y�F;t1tP�|e��Y�F ;x1tP�je��Y�v$;5|1tV�Xe��Y^]�����������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U���S�u�M��k���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�2����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M���j���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�1N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��1��+�1;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�1N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���1A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�1��1��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硠1��1�3�@�   ��1�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�1��M���Ɂ�   �ً�1]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�1N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��1��+�1;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�1N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���1A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�1��1��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硸1��1�3�@�   ��1�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�1��M���Ɂ�   �ً�1]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�@#3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u�Z���SSSSS�    葻����3��N  �U�U��< t<	t<
t<uB��0�B���/  �$���Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�q#  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  �5��`�E�;���  }�عp6�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[��R���Ðա)������/�C������������U���t�@#3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uhD�Qf��t��   �u��u;h<�;�u0��u,h4�CjP������3���tVVVVV褲�����C�*h,�CjP������3���tVVVVV�x������C3��q  �ʋ�i�M  �������Ck�M��������3���f�M�5�ۃ�`�E�f�U�u�}�M�����  }�p6�ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��I���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95�S��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��?���Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ��U��j
j �u�Q  ��]���U��SVWUj j h���u�z   ]_^[��]ËL$�A   �   t2�D$�H�3��,D��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    �@#3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ��1�SQ��1�L$�K�C�kUQPXY]Y[� ����������������Q�L$+ȃ����Y�*  Q�L$+ȃ����Y�  ��U��QQ�EV�u�E��EWV�E��  ���Y;�u�|��� 	   �ǋ��J�u�M�Q�u�P����E�;�u����t	P�|��Y�ϋ������S�����D0� ��E��U�_^��jhp�Wi������u܉u��E���u�U|���  �:|��� 	   �Ƌ���   3�;�|;�Sr!�+|���8�|��� 	   WWWWW�H������ȋ������S��������L1��u&��{���8��{��� 	   WWWWW������������[P�  Y�}���D0t�u�u�u�u�������E܉U���{��� 	   �{���8�M���M���E������   �E܋U��h����u�@  YË�U���  �g  �@#3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�{���0��z��VVVVV�    �5���������  SW�}�����4��S�����ǊX$�����(�����'�����t��u0�M����u&�z��3��0�z��VVVVV�    �ʢ�����C  �@ tjj j �u�~������u�i  Y����  ��D���  �V���@l3�9H�������P��4�� ���������`  3�9� ���t���P  �����4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�J���Y��t:��4���+�M3�@;���  j��@���SP�[  �������  C��D����jS��@���P�7  �������  3�PPj�M�Qj��@���QP�����C��D����h������\  j ��<���PV�E�P��(���� �4������)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�������  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@����D  Yf;�@����h  ��8����� ��� t)jXP��@����  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4������B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4������b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �h���;���   j ��,���P��+�P��5����P��(���� �4�����t�,���;�������@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�����t��,�����@��� ��8��������@�����8��� ul��@��� t-j^9�@���u�t��� 	   �t���0�?��@����t��Y�1��(�����D@t��4����8u3��$�Ft���    �Nt���  ������8���+�0���_[�M�3�^�-:����jh��a���E���u�t���  ��s��� 	   ����   3�;�|;�Sr!��s���8��s��� 	   WWWWW�������ɋ������S��������L1��t�P��  Y�}���D0t�u�u�u�.������E���ls��� 	   �ts���8�M���E������	   �E��`����u�1  YË�U����Bh   �R��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u��r��� 	   3�]�V3�;�|;�Sr��r��VVVVV� 	   �������3���ȃ������S���D��@^]ø�1á�SVj^��u�   �;�}�ƣ�SjP�5R��YY�hC��ujV�5�S�R��YY�hC��ujX^�3ҹ�1��hC��� ����`4|�j�^3ҹ�1W�������S����������t;�t��u�1�� B��P2|�_3�^��  �=9 t��  �5hC�?7��YË�U��V�u��1;�r"��@4w��+�����Q�Uf���N �  Y�
�� V���^]Ë�U��E��}��P�(f���E�H �  Y]ËE�� P���]Ë�U��E��1;�r=@4w�`���+�����P�e��Y]Ã� P���]Ë�U��M���E}�`�����Q��d��Y]Ã� P���]Ë�U��EV3�;�u��p��VVVVV�    ������������@^]á@#��3�9�B����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�Pp��j^SSSSS�0舘�������V�u�M��<���E�9X��   f�E��   f;�v6;�t;�vWSV�5������o��� *   ��o��� 8]�t�M��ap�_^[��;�t2;�w,��o��j"^SSSSS�0�
�����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�h�;�t9]�^����M;�t�������z�D���;��g���;��_���WSV�94�����O�����U��j �u�u�u�u�|�����]Ë�U����@#3ŉE�j�E�Ph  �u�E� �����u����
�E�P�\���Y�M�3���4���Ë�U���4�@#3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5���M�QP�֋����t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��4�����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�"2��Y;�t	� ��  ���E���}�9}�t؍6PW�u���2����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�h���t`�]��[�h�9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�1M��YY�E�;�t+WWVPV�u�W�u��;�u�u���2��Y�}���}��t�MЉ�u�茬��Y�E��e�_^[�M�3��!3���Ë�U����@#3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�S1���Ë�U���VW�u�M��7���E�u3�;�t�0;�u,�k��WWWWW�    �I������}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�����M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&�qi���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9�Auh@/�P������]����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��MS3�;�VW|[;�SsS������<��S�������@t5�8�t0�=�8u+�tItIuSj��Sj��Sj�������3���9h��� 	   �Ah������_^[]Ë�U��E���u�%h���  �
h��� 	   ���]�V3�;�|";�Ss�ȃ������S����@u$��g���0��g��VVVVV� 	   ����������� ^]�jh��T���}����������4��S�E�   3�9^u6j
�<\��Y�]�9^uh�  �FP� ���YY��u�]��F�E������0   9]�t�����������S�D8P����E��`T���3ۋ}j
��Z��YË�U��E�ȃ������S���DP���]Ë�U����@#3ŉE�V3�95�7tO�=D8�u�g  �D8���u���  �pV�M�Qj�MQP����ug�=�7u�����xuω5�7VVj�E�Pj�EPV��P�h��D8���t�V�U�RP�E�PQ� ���t�f�E�M�3�^�B,������7   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��]2���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�7���YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p������E�u�M;��   r 8^t���   8]��e����M��ap��Y����Ke��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p������:���뺋�U��j �u�u�u�������]�jh���Q��3ۉ]�j�Y��Y�]�j_�}�;=�S}W�����hC�9tD� �@�tP�  Y���t�E��|(�hC��� P�T��hC�4� *��Y�hC�G��E������	   �E��Q���j�@X��YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�C���YP�������;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�����P�  Y��Y��3�^]�jh��P��3��}�}�j�MX��Y�}�3��u�;5�S��   �hC��98t^� �@�tVPV�����YY3�B�U��hC���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�hC�4�V�����YY��E������   �}�E�t�E��P���j�V��Y�j����Y����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h����D8áD8V�5����t���tP�֡@8���t���tP��^Ë�U��SV�uW3����;�u��a��WWWWW�    �&�������B�F�t7V�{���V����  V�����P�   ����}�����F;�t
P�$'��Y�~�~��_^[]�jh�N���M��3��u3�;���;�u�la���    WWWWW裉���������F@t�~�E��N���V����Y�}�V�*���Y�E��E������   �ՋuV�����Y�jh8�N���E���u��`��� 	   ����   3�;�|;�Sr��`��� 	   SSSSS�������Ћ����<��S��������L��t�P�����Y�]���Dt1�u�g���YP����u���E���]�9]�t�z`���M��]`��� 	   �M���E������	   �E��M����u�)���YË�U��V�uWV� ���Y���tP��S��u	���   u��u�@Dtj�����j�������YY;�tV�����YP����u
�����3�V�����������S����Y�D0 ��tW��_��Y����3�_^]�jhX�L���E���u�_���  �w_��� 	   ����   3�;�|;�Sr!�i_���8�O_��� 	   WWWWW膇�����ɋ������S��������L1��t�P�g���Y�}���D0t�u�����Y�E����^��� 	   �M���E������	   �E��L����u�����YË�U��V�u�F��t�t�v�4$���f����3�Y��F�F^]�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%��������������h@��T!��Y����̃=h8 uK�`8��t�p8�Q<P�B�Ѓ��`8    �l8��tV����r��V蚜�����l8    ^�                                                                                                           � � � � �   . B P \ j t � � � � � � � �  $ : T l � � � � � � � 
   : F b � � � � � � �   " , 8 J V f � � � � � � �   . @ P ` v � � �         0�        !��6�;�X\�        ���                    ��M       {   @ @� bad allocation            �?        � � `   Render Elements Thread      7�A`���?<@2  �� �� @
@�P��� About Render Elements   Help    Mental Ray Camera Tags  VRay Camera Dome Tags   VRay Physical Camera Tags   VRay Compositing Tags   Sketch Style Tags   Sketch Render Tags  Compositing Tags    Materials   Active Camera   Render Settings Layers  Objects Save As Default Preferences Options Clean Material Editor   Delete All Elements Delete Checked Elements Set Render Camera on Checked Elements   Set Selected Layers on Checked Elements Set Selected Tags on Checked Elements   Set Selected Objects on Checked Elements    Update Checked Elements Invert Checked Elements Uncheck All Elements    Check All Elements  Edit    to  Change Frame Range      As Save Project (One Tex Folder)    As Save Project As Save File (Into Folders) As Save File    Generate .C4D Files Generate Preview Image  Record Element  Rename  Delete  Load    res default_image.tif   myBitmapButton  Render Elements tif Bitmap  You must select a camera!   (p2 t �n@n�n t pn`n/       :   0       *       �OA_RE An error has occurred while saving the Render Element!  Could not create directory to save Render Element    in!    c4d Illum   gi  illum   icon.tif        c:\program files\maxon\r12final\plugins\renderelements_0_7_13\source\renderelements.cpp tex Render Elements V   .  (c) 2011 Adam Swaab. pdf help    RE_Manual   Delete Bitmap Preview Folder     ?  You must check at least one render element! Choose a Directory to Save Generated Files      Warning! This will overwrite files in the chosen directory if they have the same name as your selected Render Elements! Are you sure you want to delete this element?  This cannot be undone.   You must save your document before you can generate preview images. Render Elements - Generating Preview Image  Render Elements - Saving Date and Time  Render Elements - Saving Layer Settings Render Elements - Saving Camera Settings    Render Elements - Saving Object and Tag Settings    Render Elements - Saving Render Settings        An element with that name already exists.  Do you want to overwrite it? You must enter a name for this element. Error! New RE Directory could not be created!   A Render Element directory with the same name already exists in that location.  Should I overwrite it?  �8��������5Ћ�0�@� �p�������P�`�P�������`�p�����Џ����    c:\program files\maxon\r12final\plugins\renderelements_0_7_13\source\renderelementsnode.cpp Render Elements Node    c:\program files\maxon\r12final\resource\_api\c4d_resource.cpp  #   M_EDITOR    c:\program files\maxon\r12final\resource\_api\c4d_file.cpp  @�p� ����c:\program files\maxon\r12final\resource\_api\c4d_general.h %s     T� ����     �f@-DT�!	@� �� � �0�@�P��`�      Y@     @�@� �� � �0�@�P��P�H�����`�p���0���P���p�c:\program files\maxon\r12final\resource\_api\c4d_gui.cpp   � �� � �0�@�P����    � �� � �0�@�P��@������ �P`@Progress Thread 0%  ~   %       ����MbP?`pc�H�Pc    c:\program files\maxon\r12final\resource\_api\c4d_baseobject.cpp    � n    c:\program files\maxon\r12final\resource\_api\c4d_basebitmap.cpp    c:\program files\maxon\r12final\resource\_api\c4d_basetime.cpp            �? �Ngm��C   ����A  4&�k�  4&�kCc:\program files\maxon\r12final\resource\_api\c4d_pmain.cpp     �������������c:\program files\maxon\r12final\resource\_api\c4d_libs\lib_ngon.cpp  �    c:\program files\maxon\r12final\resource\_api\c4d_gv\ge_mtools.cpp  PP���������a a ,��                      �?      �?3      3            �      0C       �       ��              e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    �>?          �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow         �������             ��      �@      �              �?5�h!���>@�������             ��      �@      �            	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        � ���������������������������������������������|�p�l���h�d�`�\�X�T����P�L�H�D�@�<��8�4�0�,�(�$� ������������������������`�@� � �������|�T�8�(�$���������������`�8����������T�(����GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           @#�   RSDS�c�R
O�ո��r�   C:\Program Files\MAXON\R12Final\plugins\RenderElements_0_7_13\obj\RenderElements_Win32_Release.pdb               �           ��            ����    @   �          ����    @   $           4                8 P           `l�    8        ����    @   PP         ����    @   �           ��               ���    h        ����    @   ��         ����    @               �                � <           L\��    �        ����    @   <           ���    �        ����    @   x           ����    �        ����    @   �            �             $���    �        ����    @                  $            0!h           x�    0!        ����    @   h            L!�           ���    L!       ����    @   �            P �            p!            ,�    p!       ����    @               �!\           lt    �!        ����    @   \            �!�           ���    �!       ����    @   �            �!�            ��    �!       ����    @   �           <D    �!        ����    @   ,            "t           ��    "        ����    @   t            $"�           ��D    $"       ����    @   �            �             �"           ,4    �"        ����    @               �"d           t|    �"        ����    @   d            �"�           ��D    �"       ����    @   �            �"�               �"        ����    @   �            #@           PX    #        ����    @   @            @" �h ��                     ����    ����    ����!�2�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    �����    �����    ����    ����    `����    l����    ����    ����    �    ����    ����    ������    ����    ����    ����    �$    ����    ����    ����    �)    ����    ����    ����h6�6    ����    ����    ����    �T    ����    ����    ����    yX    ����    ����    ����    �[    ����    ����    ����    �j    ����    ����    ����    l    ����    ����    �����mn    ����    ����    ����MnQn    ����    ����    ����    Gp    ����    ����    �����p�p    ����    ����    ����D�`�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �        ������    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��         �  �                     � � � � �   . B P \ j t � � � � � � � �  $ : T l � � � � � � � 
   : F b � � � � � � �   " , 8 J V f � � � � � � �   . @ P ` v � � �     �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �GetLastError  �HeapFree   GetProcAddress  �GetModuleHandleA  �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �InterlockedIncrement  �SetLastError  �InterlockedDecrement  !Sleep ExitProcess �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA � DeleteCriticalSection �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW zWideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  >UnhandledExceptionFilter  SetUnhandledExceptionFilter �WriteFile �LeaveCriticalSection  � EnterCriticalSection  TVirtualAlloc  �HeapReAlloc -TerminateProcess  �GetCurrentProcess �IsDebuggerPresent [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �RtlUnwind �LoadLibraryA  �InitializeCriticalSectionAndSpinCount �GetLocaleInfoA  ZRaiseException  �LCMapStringA  MultiByteToWideChar �LCMapStringW  =GetStringTypeA  @GetStringTypeW  �SetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW x CreateFileA C CloseHandle AFlushFileBuffers  KERNEL32.dll                  ��M              � �   ��    RenderElements.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   |�|�L�    .?AVREThread@@  L�    .?AVC4DThread@@ L�    .?AVREDialog@@  L�    .?AVGeDialog@@  L�    .?AVCommandData@@   L�    .?AVBaseData@@  L�    .?AVRE@@    |�L�    .?AVNodeData@@  L�    .?AVSceneHookData@@ L�    .?AVRenderElementsNode@@    |�|�|�|�|�|�|�|�|�L�    .?AVGeListView@@    L�    .?AVSimpleListView@@    |�L�    .?AVGeModalDialog@@ L�    .?AVGeUserArea@@    L�    .?AVSubDialog@@ L�    .?AViCustomGui@@    |�|�|�|�L�    .?AVGeSortAndSearch@@   L�    .?AVNeighbor@@  L�    .?AVDisjointNgonMesh@@  |�|�|�|�|�|�|�|�|�|�|�|�|�|�|�|�|�L�    .?AVGeToolNode2D@@  L�    .?AVGeToolDynArray@@    L�    .?AVGeToolDynArraySort@@    L�    .?AVGeToolList2D@@  |�|�|�u�  s�  |�L�    .?AVtype_info@@             N�@���D        fmod         t B�ABtAB�AB�A�A�A�ABB�ABsqrt    �g�g�g�g�g�g�g�g�g�g|�            ���������    �����
                                                                   x   
         (�   ��	   ��
   8�   �   ��   ��   ��   T�   ,�   ��   ��   ��   t�   �    ��!   ��"   @�x   ,�y   �z   ��   ��   ��                                                                                                                                                                                                                                                                                                                   	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 ?                     ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ���dCjCoCuCzC�C�C�C�C�C�C�C�C�C�CDD>DCD]DbD�D�D�D�D�D�DEE&E:EREfE�E�E�E�E�E�E�E
F*F/FIFNFnF�F�F�F�F�F�F�FG&G>GRGrGwG�G�G�G�G�G                                                                                                                                                                                                                                                                                                                                      abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     0)�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    �����C                                                                                              X.            X.            X.            X.            X.                              X1        �� 	�0`.   `.0)        �&         ��   ��   t�   x�   �   �!   �   l�   d�   T�   �   �   8�   4�    0�   L�   D�   �   <�   �   �   �   �   �"   �#   �$   �%   �&   |      �      ���������              �       �D        � 0     ��    ($  �
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
x
�
p
h
`
T
L
@
4
0
,
 

 
	         �0.   T1�B�B�B�B�B�B�B�B�BX1   .                 ���5      @   �  �   ����              �            �C    �C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �p     ����    PST                                                             PDT                                                             p4�4����        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
       ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                           �   E0d0u0�0�0�0�01141d1x1�1�1�1�1�1$2a2�2�233�3�3�3V4_4u4�4�4�4�4�46/6J6e6�6�6�6�6�67"7=7X7s7�7�7�7�7858P8k8�8�8�8�8�8+9�9�9':9:L:b:t:�:�:�:�:�:	;+;X;j;{;�;�;�;�;<Z<q<�<�<�<�<�<�=�=�=�=�=>>3>Q>c>t>�>�>�>�>�>?)?:?\?�?�?�?�?      `  0*0;0[0m0~0�0�0�0�0�01<1N1_11�1�1�1�122&2L2]2o2�2�2�2�2�2�23-3>3`3�3�3�3�3�34484y4�4�4�4�4�4�455&575R5d5v5�5�5�5�5�5�56 616L6^6p6�6�6�6�6�6�6�67!7<7X7j7{7�7�7�7�7�788%8@8\8n88�8�8�8�8�899$9?9Q9c9t9�9�9�9�9�9�9::/:A:S:d:�:�:�:�:�:�:�:;;1;C;T;p;�;�;�;�;�;�;�;<!<3<D<`<r<�<�<�<�<�<�<==(=9=U=g=x=�=�=P>`>�>�>�>?F?n?�?�?�?   0  �   060^0�0�0�0�01.1N1n1�1�1�1�12E2e2�2�2�2�23%3E3e3�3�4�4h5�5�526H6j6�6�6�677:7P7q7�7�7�728B8�8�8�89919�9�9�9�9$:A:Y:�:�:I;d;�;�;�;<5<�<�<�<
=:=I=i=�=�=�=�=>'>W>f>�>�>�>�>?$?D?�?�?�?   @  �   0&0N0l0�0�0�0�0181`1~1�1�1�12)2D2l2�2�2�2�23>3\3�3�3�3�34.4V4t4�4�4�4 5(5F5n5�5�5�5�56@6^6�6�6�6�67*7R7p7�7�7�7�7808X8v8�8�8�89*9H9p9�9�9�9�9:B:`:�:�:�:�:;2;Z;x;�;�;�;<,<J<r<�<�<�<�<=D=b=�=�=H>r>�>�>�>?;?Y?w?�?�?�? P    
0/0�0�0_1v1�1�1�1�1�1	2"2;2T2m2�2�2�2<3R3w3�3�3�3�34"4C4W4u4�4�4�4�4�45<5P5n5�5�5�5�5�5656K6k6�6�6�6�6�6787N7n7�7�7�7�7�78;8O8m8�8�8�8�8�8949H9f9�9�9�9�9�9:-:A:_:�:�:�:�:�:;&;:;X;y;�;�;�;�;�;<3<Q<r<�<�<�<�<�<=,=J=k==�=�=�=�=>%>C>d>x>�>�>�>�>
??<?]?q?�?�?�?�? `  �   0050V0j0�0�0�0@1�1�102�2�2 3p3�3�34F4\4z4�4�4�4�4�45<5`5�5�5�5 66!6H6�6�6�6�6�6A7Q78%8N8�8�8�89:9S9x9�9�9�9:�:�:�:�:;2;|;�;<8<]<�<�<�<�<=g=�=�=�=�=c>�>�>�>�>�>�?�?�? p  �   	0B0Z0�0�0�0�0u1�1�1�1�12;2�23&3B3Y3r3�3�3�3D4r4�4�4�4�4�45525P5j5�5�5�56'696^6p6�6�6�6�6�6�67+7H7�7�7�7888G8�8�89>9p9�9�9�9�9�9:0:H:z:�:;=;O;f;�;�;�;�;<N<x<�<�<�<�<'=?=V=z=�=�=�=>)>[>�>�>�>�>
?4?L?c?�?�?�?�? �     040�0�0�0�0�01/1I1e1�1�12272Q2�2�2�2�2�3�3�3�3�34-4E4]4u4�4�4�4a5s5�5�5�5�5�56\6k6�6�6�6 77&7;7P7d7�7�7�7	8!8@8R8p8�8�8�8�8939V9w9�9�9�9�9�9:0:W:h::�:�:�:�:;!;C;V;j;�;�;�;�;"<F<b<�<�<�<�<�<==4=M=f==�=�= >>F>t>�>�>?-?N?s?�?�?�?�?�?�? �    0!0:0Y0�0�0�01161U1g1�1�1�1�12 2C2y2�2�2�2�2333�3�3�3�3424^4s4�4�4�4�4�4"535h5x5�5�5�566+6H6�6�6�6�6�6	7#7=7W7q7�7�7�7�7818R8i8�8�8�8�8�89(9?9[9y9�9�9�9�9::-:D:d:�:�:�:.;=;k;�;�;�;�;�;<<)<F<`<u<�<�<�<==E=b=�=�=�=�=�=�=>(>A>Z>s>�>�>�>�>0?I?a?y?�?�?�?�?�?   �  ,  0"0v0�0�0�0�0121X1j1~1�1�1�1�1�1'2�2�2�23V3�3�3�3�3�34$464q4�4�4�4�4�4	5'5N5p5�5�5�5"636X6j6�6�6�6�6�6�67	7"7D7b7�7�7�7�7�78'8:8N8`8r8�8�8�8�8�89B9W9�9�9�9�9�9�9:":4:[:m:�:�:�:�:�:�:;;);:;O;d;�;�;�;�;�;�;<%<N<e<z<�<�<�<�<�<:=O=x=�=�=�=�=�=>&>;>e>z>�>�>�>�>�>?#?;?W?q?�?�?�?�?�?   �  \  0.0>0`0v0�0�0�0�0�0(1=1E1j1y1�1�12-2`2�2�2�23:3P3c3v3�3�3�3�3�3�34)414G4^4s4�4�4�4�4�45515I5c5x5�5�5�5�5�5�56#676L6g6~6�6�6�6�6�67)7?7_7t7�7�7�7�7�7�7�78/8N8j8~8�8�8�8�8�89(9=9F9]9r9�9�9�9�9�9::2:G:_:s:�:�:�:�:�:�:�:�:
;";+;@;\;s;�;�;�;�;�;<(<?<^<s<�<�<�<�<�<='=<=W=n=�=�=�=�=�=>>.>J>_>t>�>�>�>�>�>�>??.???Q?Z?r?�?�?�?�?�? �  �   0#080L0a0s02C2n2�2�2�2\3�3�3�3�3�3�3	44/4E4Y4r4�4�4�4�455.5B5]5�5�5�5�5�5V6m6�6�6�6�67I7e7�7�7 888/8C8\8�8�8�8@9Q9c9z9�9�9):E:Z:l:�:�:�:�:�:�:;;M;];y;�;�;<%<W<|<�<�<�<�<�<='=>=]=r=�=�=�=>>/>�>�>�>�>7?�?�?�?�?   �  �   0�0�0�01)1>1U1t1�1�1�1�1�12%2P2�2�2�23�3�3�3�3�34#4:4Y4n4�4�4�455.5C5U5f5�5�5�5	66X6m6�6�6�6�67/7�7818F8X8l8~8�8�8�8�8�8999I9e9�9�9�9:C:h:�:�:�:;5;x;�;%<:<N<i<=1=F=a=x=�=�=�=�=�=
>9>N>b>w>�>? ?5?P?�?�? �  �   0$0@0U0k0�0�0�0�0�051J1_1s1�1�1�1�122<2S2r2�233Q3s3�3�3�3�3�344 414C4L4^4p4�4�4�4
55'6G6V6n6�6�6�6�6�6�6F7r7�7�7�7�78T8�8�8�8�8�8�9 :A:S:e:y:�:�:�:�:�:
;;3;Q;e;w;�;�;�;�;�;<<.<C<q<�<f=�=�=�=>�?   �  �   030v0�0�0�0�0�0�011-1S1g1�1�1�1�1/2T2u2�2�2�223X3k3�3�3(4]4r4�4�4^5s5�5�5�5�5�56686O6{6�6�6�6�6K7`7u7�7�7�7?8f8{8�8�8�8�8�89909G9v9�9�9�9::*:H:�:�:�:�:;�;<�<�<�<�<C=?W?v?�?�?�?�?�?�?�?   �   040H0~0�0�0�0151V1�1�1�1282K2i2�23K3`3u3�3L4a4v4�4�4�4�4�45&5=5i5~5�5�5�586M6b6}6�6�6&7N7c7w7�7�7�7�7�78'8>8�8�8�8�8�8�89%9i99�9�9�9s:�:;>;S;�;�;�<�<�<�<�<�<�<(=�=�=�=>>9>T>o>�>�>�>�>�>?(?g?~?�?�?  �   0?0V0{0�0�0�01D1j1�1�1�1�1�1�1252P2l2�2�2�2�2
3"3<3X3v3�3�3�3�3�3�3#4:4�45�5�5�5�5�5%6N7`7r7z7�7�7�7�7�7:8K8]8f8�8�899J9\9e9}9�9�9�9�9 :7:N:h:�:�;�;�;�;�;<=(=f=�=�=>I>�>�>"?8?J?�?     �   #090W0m00�0�0�0�01+1=1Q1p1�1�1!2E2Z2�2�2�2 33-3�3�3�344(4<4E5f5�5�5�5�5�56#6>6Y6t6�6�6.7M7�7�78%8�8�8�8�9�9�9R:m:�:;:;Y;�;<&<�<�<�<�=�=�=S>n>�> ?;?Z?�? 0    0'0z0�0�0�0R1a1�1�1�1�1�1�2�2�2�23[3n3�3�3�3�3�3�3�5�5)6T6i6�657F7�7�7�7�7�7B8I8f8�8�8�89K9�9�9�9�9�9�9:!:.:F:Y:k:}:�:�:�:�:�:;;4;E;X;�;�;�;�;�;�;�;�;<&<D<V<r<�<�<�<�<�<�<=&=B=S=f=�=�=�=�=�=�=�=>>6>T>f>�>�>�>�>�>�>�> ?6?R?d?v??�?�?�?�?   @ $  $020?0W0i0{0�0�0�0�0�0�01(1D1V1h1q1�1�1�1�1�122-2N2d2�2�2�2�2�2�2373d3�3�344$464@4[4w4�4�4�4�45-5V5x5�566(616D6�6�6�6�677,7R7o7�7�7T8i8�8�8'949a9r9�9�9�9�9�9�9:%:3:Q:b:�:�:�:�:�:;,;@;P;t;�;�;�;�;�;�;<,<@<O<_<p<�<�<�<�<=$=D=d=�=�=�=�=�=>4>T>�>�>�>�>�>!?4?d?�?�?�?�?�?   P   010A0Q0d0�0�0�0�01$1D1d1�1�1�1�12252'3X3j33�3�3�3D4o4�4�4�45$5D5d5�5�5�5�56!646d6�6�6�6�6�677-7;7J7\7�7�7�7�7�78$8Q8a8q8�8�8�8�8�8�8�899,9T9t9�9�9�9�9:4:T:t:�:�:�:�:;);E;];w;�;�;�;�;<4<T<t<�<�<�<�<�<�<="=1=A=S=t=�=�=�=�=�=>">7>Q>b>�>�>�>�>�>�>1?D?t?�?�?�?�?�? `    0$0D0d0�0�0�0�01$1D1d1�1�1�1�12$2D2d2�2�2�2 3$3D3d3�3�3�3�34$4D4d4�4�4�4�45$5D5d5�5�5�5�56$6D6a6t6�6�6�6�67!717A7T7t7�7�7�7�78$8I8j8�8�8�8�9�9::-:`:u:�:�:;4;Q;d;�;�;�;�;<D<t<�<�<�<�<E=Q=[=a=f=�=�=�=�=>1>D>a>t>�>�>�>??#?(?T?k?�?�?�?   p �   !0A0a0�0�0�01<1d1�1�12%2�2�2	3%3�3�3	4,4H4l4�4�4�4�4M5e5�5<6a6�6�67$7D7d7q7�7�7�78$8A8T8�8�8�8�89/9O9b9�9�9�9�9:T:t:�:�:�:�:$;D;t;�;�;�;<4<q<�<�<�<�<=4=T=t=�=�=�=�=>$>D>d>�>�>?#?�?�? � �   !0G0�01:1]1�1�12�2�2�2>3^3s3�34D4q4�4�4�5�5�5S6|6�6#7L7t7�78#8�8979�9�9:7:�:�:;|;�;<D<�<�<�<n=�=�=�=Q>�>,?T?t?�?�?�?�?   � �   00@0d0�0�0�0141T1t1�1�1�12B2`2�2�2�2�2
3G3V3�3�3�3�3444�4�4�4�4�4!5D5t5�5�5�5�56D6t6�6�6�6�6�67W7�7�7�7'8b8�8�8�8$9A9T9�9�9�9�9:4:T:�:�:�:;4;d;�;�;�;�;<4<T<t<�<�<�<�<�<==4=T=t=�=�=�=�=4>T>t>�>�>�>�>�>?$?D?d?�?�?�?�? � �   040T0t0�0�0�0�0111D1d1�1�12$2D2d2�2�2�2�23$3D3d3�3�3$4S4�4�4$5Q5t5�5�5�5646T6q6�6�6�6�6�6747i7}7�7�7888d8�8�8�899&9T9r9�9�9�9�9:$:D:d:�:�:�:�:;";D;j;�;�;�;�;�;<"<2<T<n<�<�<�<�<�<=D=\=�=�=�=�=�=>,>U>�>�>�>�>�>?;?N?�?�?�?�? � �   $0D0d0�0�0�0�0141T1q1�1�1�1�1242T2t2�2�2�2�2343T3q3�3�3�3�3�34!4D4Y4k4�4�4�4�4�4�4�4�5�5�5646d6�6�67(7U7a7u7{7�7�7�7�78D8q8�8�8949d9�9�9�9 :�:�: ;6;d;�;�;�<�<�<�<�<=4=a=�=�=�='>@>�>�>�>:?\?�?�?�? � �   0,0{0�0�0D1�1�1�182Q2l2�2�2�2�2�2'393�3�3�3�3 44V4�4�4�4�45>5U5{5�5�5�56)6V6h6�6U7]7�78[8�8�8'9]9�9�9:0:i:�:�:�:6;k;�;�;<1<N<t<�<4=�=>E>�>�>�>?]?�?�?   � x   20�0�0�01R1�1�1�1�122Q2�2�2�2�3�3#4�4�45`5�56s6�6$7s7�738�8�8S9�9:s:�:0;�;�;C<�<===�=>`>�>�>�> ?P?�?�?�? � �    0m0�0�0�0141n1�1�1*2{2�23^3�3�34B4d4�4�45D5�5�5�556U6n6�6�6e7j7u7�7�7�788T8�8`9�98:<:@:D:H:L:P:T:X:�:9;�;�;�;�;�;�;�;�;�;V<x<�<�<�<�<�<!=A=a=�=�=�=�=$>D>d>�>�>?D?d?�?�?   � �   00�0�0�0!1D1t1�1�12)2F2X2j2�2�2�2�2�2�2303A3U3s3�3�3�3�3�3�3444�4�4�4�4$5d5�5 646t6�6�6747t7�7�7�7�8�8959N9u9�9(:?:X:r:G;�;�;<<%<:<X<b<�<�<$=D=d=�=�=�=�=�=s>�>E?�?�?�?   �   $0T0�0�0c1�1�1�12!2a2v2�2�2�2�243q3�3�3�3�3�34D4t4q5�5�5�56"656U6�6�6�6�677Z7~7�7�78/8A8R8y8�8�8�8 99'949_99�9�9�9:>:p:�:�:8;�;�;<D<s<�<�<�<=R=�=�=�=>">;>M>i>w>�>�>�>�>
??$?7?O?d??�?�?�?�?�?�?    �   0 2�2�243�3�3Y4�4�4T5u5�56�6�6h7�748M8v8�8�8�8�8�8999V9�9�9::0:<::�:�:�:�:;.;];k;{;�<�<+=5=�=�=�=>!>A>e>�>	?�?�?   �   0U0�0�0�1�1252u2�2�253�3�3�34E4�4�45e5�5�56E6�6�6"7U7�7�78E8�8�8�8%9u9�9:E:�:�:�:;$;4;U;�;�;%<b<�<�<5=�=�=�=!>I>S>�>�>�>�>�>%?I?�?�?�?   0 �   0e0�0�0�01F1o1�1�1282v2�23!3D3�3�344t4�4�4�4�4545T5t5�5�5�5646T6�6�6�6�6!7D7q7�7�7�78A8d8�8�8�8919Q9q9�9�9�9�9:1:Q:q:�:�:�:�:;4;d;�;�;�;�;!<D<a<�<�<�<=$=T=�=�=�=>b>�>�>�>�>?4?a?�?�?�?�?   @ �   040d0�0�0�01$1D1d1�1�1�1�1212@2d2�2$3Q3d3�3�3�3414Q4�4�4�4�4515T5�5�5�56D6t6�6�67J7�7�7�78!8D8t8�8�8�8�8�89Z9t9�9�9:::�:�:�:�;�;1<E<Z<}<�<�<�<3=V==�=�=>$>h>�> ?d?t?�?�?�?   P �   )0S0g0�0�0�0�0141d1�1�1�1�1242�2�2�2�2!3A3d3�3�3�3�3D4�4�4�4�45_5~5�5�566H6c6�6�6�6�67,7F7v7�7�7�7�78?8S8h8�8�8�8919K9k9�9�9W:j:�:�:�:�:!;l;{=   ` �   *0C0�0�0�0�0'1d114383<3@3{3�3�34444T4t4�4�4�4�45515A5T5q5�5�5�5�56(6A6d6�6�6�6�6747T7t7�7�7�7818A8T8t8�8�8�8�8919O9t9�9�9�9:5:M:\:�:�:�:�:�:;;-;t;�;�;�;$<4<a<�<�<�<�<�<=A=T=t=�=�=�=�=>t>b?i?p?w?~?�?�?�?�?�? p �   0�0E1�1�1�1�1242T2q2�2�2�23$3D3d3�3�3�3�3!4�4�4!545a5�5�5�5�5636F6q6�6�6�67$7T7�7�7�7�78T8�8�8�8�8$9D9a9�9�9�9�9:4:f:{:�:!;4;d;�;�;�;�=�=�=�=�>�> � �   X0�0�0�01$1Q1a1q1�1�1�1�12D2d2�2�2�2�2�2343Q3d3�3�3�4�4:5?5�5s6�6�637F7V7�788�8�8�8�8i9�9::1:::M:�:�:�:�::;J;�<�<�<{= >>>>>#>*>1>8>?>F>M>T>[>b>i>p>   � �   $0.080B0L0V0`0j0t0~0�0t1�1�1�1�1!2d2�2�2�2�2�23343N3�3�3�3�3�3�3�3�3�3�45B5u5�5E6�6�67U7�7�728b8�8�859u9�9�9R:�:�:2;b;�;�;<2<e<�<=8=L=\=z=�=�=%>u>�>?U?�?�?   � t   E0�0�0"1b1�1�122x2�223x3�324u4�45e5�56R6�67�78U8�8�89e9�9:E:�:�:5;�;�;<e<�<=e=�=�=>->e>�>�>5?�?�?   � D   %0u0�0%1�1�12U2�2�2%3e3�34^4�4�45]5�5�5,66�6|7�7�78�8�8 � ,   2Q<q<�<�<=U=�=�=%>b>�>�>?B?u?�?�? � l   50r0�0�0121e1�1�152�2�23E3�3�354�4x6�6.9�9�9�9�9�9�:�:�:�:R;`;�;�;N<\<�<�<�<�<�=�=>!>�>�>�>�>�?�? � X   �3=4M4|5�56D6K6f6�6�6�67]7�7�7�8�8�9:S:�:�:�:�:d<�<$=>$>D>t>�>�>?4?d?�?�?�? �    0}0�0�01111 1'1.181B1I1P1W1^1e1l1s1z1�1�1�1�1�1�1)2�2U3f4k4q4u4{44�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4Q5V5`5�5�5�5�5 66!6Q6m6�6�67r7}7�7898>8U8�8�8�849:9Z9�9�9:m::�:�:�:�:;Z;s;�;<<"<B<^<=O=h=o=w=|=�=�=�=�=�=�=�= >>>>>>^>d>h>l>p>�>�>�>????1?[?�?�?�?�?�?�?�?�?�?�?   �    0000a0k0x0�0�021=1O1�1�1�1�1n4�45e: ;�<==G=M=V=]=r=�=�=p>v>�>�>�>�>�>�>�>�>�>??$?8???W?c?i?u?�?�?�?�?�?�?�?�?�?�?�?�?    T  
000A0V0|0�0�0�0�01&1L1�1�1�1+2322�2�2�2�2�2�2�2�2�2�2333 3'3-343:3B3I3N3V3_3k3p3u3{33�3�3�3�3�3�3�3�3�3�3�3�3�344484>4Z4�4�4�4�4�4�4'505<5`5i5�5�5�5�5�5�5H6P6c6n6s6�6�6�6�6�6�6�6�6�6�677\7i7�7�7�7�7�7R8_8h8|8�8�8�8,949t9~9�9�9 :0:B:�:�:�:�:�:	;;P;Z;�;�;�;�;�;�=�=�=�=�=�=$>*>@>K>b>n>{>�>�>??M?f?u?z?�?�?�?�?�?�?�?     �   000(040=0E0O0U0[0}0�0�011�12R2,343L3d3�3�3�3444!4-4Q4Y4e4�4�4�455?566%676T6�6�6�6�6�6�6�6+707X7}7�7�7�7�78*878>8H8r8�8�8�8�8�8�8�8�8�8#9�9�9�9�9.<<<B<\<a<p<y<�<�<�<�<�<�<�<�<�<�<�<	====&=-=A=H=N=\=c=h=q=~=�=�=�=�=�=+>   0 �   �1�12,2f2�2~4�4�4�4�4�4575D5N67�7�7�7�7�78888 8'8.858=8E8M8Y8b8g8m8w8�8�8�8�8�8�8�8�8�8�899%9�9�9�9�9:":.:::_:h:q:~:�:�:�:�:�:�:�:�:�:;;;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;<>A>�>Q?a?m??�?�?   @ <   �0 1�12h2�2�2�2�283`3e:�;�;<�<�<�<=a>|>�>q?{?�?   P �   k0l1|1�1�1�1�1O2�2�24'4a4n4x4�4�4�4�4�4�4�455<5s5�5�5+6H6�6�67�7�7�7�7�7�7�78888A8G8P8U8d8�8�8�8�8�9�9":n:�:;k;�;�;�;�;<�<�<�<==3=�=�=�>?�?   ` �   �0�0�0�0�0�0 11-1S1q1x1|1�1�1�1�1�1�1�1�1�1�1�1V2a2|2�2�2�2�2�2�23333 3$3(3,303z3�3�3�3�3X6i8u8�9�9::a:g:s:�:�:3;�;�;�;�;<B<v<|<�<�<x=}=�=�=�=�=0>g>r>�>�>�>�>�>�>�>#?(?m?r?y?~?�?�?�?   p d   00�0�0�0�0�0�1�1�1�1�1�1�1�1�1�1�1222$2.2<2|2�2�24%4+4s5z5�6'7E7k7�7�7�7D;4<�=�=>�?   � `   �1�1�1�122	222B4�5�5�5�5�5b6k7�78q8�8�:�:�:;';5;e;�;�<�<�<�<�<===I=y=>�>�>a?   � \   20�0�0�0�0�0�01	191�1G2T4f4x4�4�4�4�4�4�45/7%8-8�8�9[:a:;	;;�;�;s<i=q=$>?�?�?   � @   G0M0]0�01D1�1�4�488888888#8'8+8/8<89/9>9j9�9�9 � <   �3�6�6	7�7�7�7@8M8f8�8�8�8�9:�:�:�;�;U<�=�>�?�?�?   � �   030�0131�12D2W2]2w2�2�2�2�2�2�2�2�233"373A3g3�3�3�3�34>4I4t5�5�56.6g6t6S7b7�7�;�;N<^<y<�<�< =;=W=�=�=�=�=>>>+>I>S>\>g>|>�>�>�>�>_?�?�? � T   0%0L0Y0^0l0G1j1u1�1�1�2�2�2�2�2�2W3�3�3'4^4h4�455'5P5�5�5 717B7J7T7f7p7�7 � ,   1,1014181<1H1L1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�5�5�5�5�5�5�5�5�5�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;0<4<8<<<@<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=(>,>0>4>8>�>�>�?�?   � �   $0(0,0004080<0@0D0H0L0�7�7?? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?     �    00000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�04<8<�<�<�<�<�<�<== =0=4=H=L=\=`=d=l=�=�=�=�=�=�=�=�=�=�=�=>> >4>8>H>L>P>T>\>t>�>�>�>�>�>�>�>�>�>�>�>�>�>?????$?<?L?P?`?d?t?x?�?�?�?�?�?�?�?�?�?�?�?  �   000 0$0,0D0T0X0h0l0t0�0�0�0�0�0�0�0�0�0�0�0 1111(181<1D1\1l1p1�1�1�1�1�1�1�1�1�1�1�1 2222(2,242L2\2`2p2t2|2�2�2�2�2�2�2�2�2�2�2333(383<3L3P3X3p3�3�3�3�3484X4d4�4�4�4�4�4�45$5(5H5h5�5�5�5�5�566(6D6H6d6h6�6�6�6�67707P7p7   �   000 080P0h0�0�0�0�0�0�011111 1$1(1,101L1l1p1�1�1�1�1�1�1�1�12$2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�233333`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4.82868:8>8B8F8J8N8R8V8Z8^8b8f8j8n8r8v8z8~8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�899
999999"9&9*9X=P>�>�>�>�>�>?(?,?0?4?8?@?D?P?T?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? 0 �   0000$0,040<0D0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1P1X1\1`1d1h1l1p1t1x1|1�1�1�1�4�4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    