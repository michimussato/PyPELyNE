MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       D
� k{� k{� k{��˼�k{�9��5k{�9��}k{�9��#k{�ݔ��k{� kz�Lk{���-k{���k{���k{�Rich k{�        PE  L ߃DT        � !  �  �     ��     �                         p	         @                   �� K   � (                            � 4}  @� 8                           �i @            � �                           .text   ��     �                   `.rdata  ��  �  �  �             @  @.data   �E   �  &   �             @  �.reloc  4}   �  ~   �             @  B                                                                                                                                                                                                                                                                                                                                                                                                h`��Ѫ Y���������������������U������D� 8���V=�  v3�^��]�h<�h�   h�j���    �� ����t���1� ����
���    h<�h�   h�j�J� ����t����� ����
���    �&� ����M������    Q�@�@�С���M�j j�hh��@Q�@�С���M�Q�@�@�С���M�j j�hd��@Q�@�С���M���(�@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�ЍE�P�ߜ ����M�Q�@�@�Ѓ������V�@�@�С���M�VQ�@�@�Ѓ���H  ����M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ�$�L  ��ul����M�Q�@�@�С���M�j j�hl��@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ��L  ��ul����M�Q�@�@�С���M�j j�ht��@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ��dt  ��ul����M�Q�@�@�С���M�j j�h|��@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ��]  ��ul����M�Q�@�@�С���M�j j�h���@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ��
d  ��ul����M�Q�@�@�С���M�j j�h���@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ��Ee  ��ul����M�Q�@�@�С���M�j j�h���@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ���f  ��ul����M�Q�@�@�С���M�j j�h���@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�Ѓ�����M�Q�@�@�С���M�j j�hx��@Q�@�С���MЃ��@Q�M��@x�Ћ������E�P�I�I�у���tZ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��M���Q�M�QP��  ���kG  ����M�Q�@�@�Ѓ���C  �M�誶 ����M�jh�  �@�@4�С���M�jh�  �@�@4�С���M�jWh�  �@�@4��j�E�Ph&� 蕞 ���M�誶 ����M�Q�@�@�С���M�Q�@�@�Ѓ��   ^��]������������V�5����t���^� V�� ���5�����    ��t���:� V�� �����    ^������U������   �S8���VW=�  v	3�_^[��]ËE=�  ��  t#�� ��  Hu۹x��q� �����_^[��]Ë��   ���   ��jjP�E�虏 ���M��>� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M����@Qj�M��@8�С���M�Q�@�@�С�����M����   ���   �Ѕ���  �E��� ��	 �
��$    �I ����M����   ��?���P���   �Ћ���؋��   �ˋRx�ҋ�����E�P�I�I�ы���A�M�QV�@�Ѓ����=� �ˉE��� �    t����M�Q�@�@�Ѓ���  �Eԋ�P��p���P��� ��蚒 ��p����� ����Mԋ@�@<�Ѕ�uT����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�M�Q�@�@�С���M�Q�@�@�Ѓ� �������@V�@�С���M�VQ�@�@�Ѓ��E�P�f)  �ȃ���tL����U�RW�@�@8�С���M�Q���W�@�@8�С���u�����P��'  P�B4���   �M��	� ����M�Qj�M��@�@8�С���M�QW�M��@�@8�С���M�Q���W�@�@8�С���u�����P��'  P�B4�С���M��]�QS�@�M��@D��C�M��]��� ����M�Q�@�@�С���M�Q�@�@�Ѓ����G�M����   ���   �Ѝ�?���;����������M�Q���h�	 �@�@D�ЍM��w� ����M�Q���   ���   �Ѓ��   _^[��]�=�  �F����aa  j �S  ����R  _^�   [��]�������U���M�\M�YM�XM�M�E]����������������U���EW�f/�v
�M�E]����f/�w��E�E]��������������U���UW�f/����v(��	f/�v(��]f/�v(��	f/�v(��ef/�wf/�v�E(�� �X�P]�(ċE� �X�P]����U���E�Mf/�v
�M�E]��E�E]����������U���M�Ef/�w(��Mf/�v
�E�E]��M�E]������������U���M�Ef/�w(��Mf/�v
�E�E]��M�E]������������U���E�Mf/�v
�E�E]��M�E]����������U���E�Mf/�w(��Mf/�v
�E�E]��M�E]������������U���E�Mf/�w(��Mf/�v
�E�E]��M�E]������������U���E�M4f/�w(��M�U,f/�w(��U�]$f/�w(ӋE��H�@]��U����E�����j ����]��E��\�fT@��\��M��E���]�U���E��f/���E�$v
耇 ��]��V� ��]��U���M�\M�YM�XM�M�E]����������������U���M$�\M�U<�E�Y��XM��M,�\M�Y��XM�H�M4�\M�Y��XM�H]�������������U���E�\Ef.���E���Dz��]��E�e�u]��U���E�M�YX��Y���X��E�Y��X��M�E]�����U���E�XE�XE�Yh��E�E]�������������U���M�Ef/�v(��E�Mf/�v�M�E]�U���E�M�Y���Y8��X��E�Y��X��M�E]�����U���]W�f/����v�X�f/�v�\��% �(��Y�f/�v!�M�\M�Y��Y��XM�M�E]����(��Y�f/�v�E]�(��Y �f/�v-�U�\U����\��Y��Y��XU�U�E]��E]�������U���}��(�ef/�vf(��f(��mf/�wf(�f/�vf(��f(�f/�wf(�f(�W�f.��X�f(П�u��Y5���u���Dz	f(��  �E�f(�f/���\��u�v����\��\��^���^u�f(��M��\��Y��f.]�E�� ��}��^���X��^}��}�f(��\��^��X��^}��}�f(��\��^��}����X��^E���Dzf(��\U��9f.ܟ��Dz�U��Xh��\��f.ݟ��Dz1�U��X���\U�W�f/����v�X�f/�v�\ЋE�E���p�@��]����U���UW�f.ן��Dz �E�Uf(�f(��0�H�P]�����]f/��-��v
�X��Y��f(�(��X��Y��\�f(��e�5��f(��Xh��Y�f/��\�v�X�f/�v�\��= �f(��Y�f/�v(��\��Y��Y��X��If(��Y�f/�v(��6f(��Y �f/�v!���(��\��\��Y��Y��X��(�W�(�f/�v�X�f/�v�\�(��Y �f/�vf(��\��Y ��Y��X��W���(��Y�f/�v(��=(��Y �f/�v)���(��\��\��= ��Y��Y��X��(��= ��\%h�W�f/�v�X�f/�v�\�(��Y�f/�v#�E�\��0�Y��H�Y��X��P]�(��Y��f/�wK�-��(��Y �f/�v/����\ӋE�\��0�Y��H�Y��X��P]�(ӋE�0�H�P]�����U���MW��U�\�f.ȟ��D{�E�\��^��E�E]������������U���MW��e�\�f.ȟ��Dzf(���U,�\��^�f.ȟ��Dzf(���]$�\��^�f.ȟ��D{�E�\��^��E� �X�P]���������U���M�\M�YM�XM�M�E]����������������U���M�UE�Ef��\�f�fY��YU,fX��X� �P]������U���M���f.ʟ��Dz�E]�W�f/�r��]��]f/�s��^�(�(��
p �E�E]�U��������U$f.ӟ��Dz�E�oE� �~Ef�@��]�W�f/�r�M��1�Ef/��E�s!(��^��o �U$W�����E�f/�r�M��)�Ef/��E�s(��^��_o �U$W��E�f/�s(f(��Mf/�sf(�����^��(o f(ȋE�E��@�E���@��]������U����eW�f.��E����Dz�E��]����f(��^�f.ӟ��Dz�E�E��7f/�s1�Mf/��M�s!(�(��^��n ����e�E��E�\�f(��mn �YE��E�E��]�������������U����]W����f.��E���Dz�U�U��   f(��^�f.���Dz�E,�E��4f/�s)�U,f/��U�s�^�(���m ����]�E��E�\��m ���f(��Ye�W��]�U�e�f.؟��Dz�U��{f(��^�f.���Dz�E$�E��4f/�s)�U$f/��U�s�^�(��Hm ����]�E��E�\��(m �]f(��YM�W��U�M�f.؟��D{x���f(��^�f.���Dz�E�E��7f/�s1�Mf/��M�s!(�(��^��l ����]�E��E�\�f(��l f(��YU��E�E��@�E���@��]�������������U���E�Mf/�v
�M�E]��E�E]����������U���M4�Ef/�w(��U,�Mf/�w(��]$�Uf/�w(ӋE��H�@]��U���E�M]������U���E�YE$�E� �E�YE,�@�E�YE4�@]�������������U���Uf.�����Dz��]����f(��\E�^��\��M�E]����U���]W����f.ٟ��Dz(��f(��\E4�^�(��\��ef.���Dz(��f(��\E,�^�(��\��mf.���D{f(�(��\E$�^��\ȋE��`�X]�������������U���E�XE���f/�vW��E�E]��\��E�E]�����������U���EW��XE4���f/�v(���\��M�XM,f/�v(���\��e�Xe$f/�w(��\ڋE��H�@]�������U���U�E$�XU�XE,�]�e4�E�X��X��Yh��Yh�f/�v�oE� f�X]��oE$� f�`]���������������U���E�Mf/�v
�E�E]��M�E]����������U���E�M4f/�w(��M�U,f/�w(��U�]$f/�w(ӋE��H�@]��U�����f(�f(��\M�\E�Y��\��U�E]��U������Ef(��\Mf(��\E$�Y�f(��\�f(��\M� f(��\E,�Y�f(��\�f(��\M�@f(��\E4�Y��\��P]�������������U���E���f.����DzW��E�E]��\��E�^��E�E]���U���]W����f.ٟ��Dz(��f(��\��]4�^��ef.���Dz(��f(��\��e,�^��Ef.����D{�U$�\��^ыE��`�X]����������U���E�E]������U���E�XE$�E� �E�XE,�@�E�XE4�@]�������������U���U�E$�XU�XE,�]�e4�E�X��X��Yh��Yh�f/�v�oE� f�X]��oE$� f�`]���������������U������]f/�v
�E�M��]����f(�(��\M�\��Y��Y���\��U�E]���������������U���5���e4f/�����-��v�]�Y��Y��!f(�f(��\M�\�f(��Y��Y��\��},f/�v�e�Y��Y�� f(�f(��\M�\�(��Y��Y��\��}$f/�v �U�E�Y��`�X�Y��]ËEf(��\Mf(��\��`�X�Y��Y��\��]������U����������ef/�vC�M(��Y������\�(��Y��Y���Y��Y��X��$�$��]��E�Wr �M�Y������\��\]�Y��M�Y���Y��X��$�$��]�����U�����m4�����f/�v9�%��(�����Mf(��Y��\�(��Y��Y��Y��Y��E�E�q �%��f(��M4����E�Y��Y��\��Y�f(��\M4�Y��m,�X����f/��\$v)�M(��Y�f(��\�(��Y��Y��Y��Y��E�E�&q �%��f(��M,����E�Y��Y��\��Y�f(��\M,�Y�����X��$�]$f/�v)�M(��Y��\�(��Y��Y��Y��Y��X��A�E�p �M$�Y������\��\U$�Y��M�Y���Y��XЋE�$�@�D$��@��]������U������Uf/��]v@W�f.؟��Dz
�E�E]��Y�����(��\��^��\��M�E]����f.؟��DzW��E�E]��\��\��Y���^��U�E]���������U���-��W��U4f/��=���]�%��v(f.ٟ��Dz(��<�Y�f(��\�(��^��\��#f.ܟ��Dz(���\�f(��\��Y��^��],f/��uv(f.���Dz(��<�Y�f(��\�(��^��\��#f.����Dz(���\�f(��\��Y��^��u$f/�v9�mf.���D{L�Y�f(ċE(��\��X�P�^��\��]��Ef.ğ��D{(��\��\��Y��^̋E��X�P]����U������Ef/�v6�Y������XEf/�vW��E�E]��\��E�E]��\��Y���XE�E�E]����������U�����W��E4f/��5���-��v�Y��XEf/�v(���\���\��Y��XE�M,f/�v�Y��XMf/�v(���\���\��Y��XM�e$f/�v)�Y��Xef/�w*�E(��\��H�@�]�(��\��Y��XU�E��H�@]��������U������Ef/�v'�Y���Mf/�v
�M�E]��E�E]��\��M�Y��f/�v
�M�E]��E�E]���������U������E4f/�����]v
�Y�f/���\��Y�f/�w(��E,f/��ev
�Y�f/���\��Y�f/�w(��E$f/�v�M�Y�f/���\��M�Y�f/�w(ȋE��`�X]�����U���%��W��Mf/��m���v,f.���Dz(��?�Y��f(��\�(��^��\��"f.���D{(�\�f(��\��Y���^�f/�w
�U�E]��]�E]���U���%�����M4W�f/��-���u���v(f.���Dz(��7�Y�f(��\�(��^��\��f.���D{!�\�f(��\��Y��^�f/�w�U���]��M,f/��uv(f.���Dz(��7�Y�f(��\�(��^��\��f.���D{ �\�f(��\��Y��^�f/�wf(��f(��M$f/��uv(f.���Dz(��7�Y�f(��\�(��^��\��f.���D{�\�f(��\��Y��^�f/�v(ӋE�E���x�@��]���������U���E�\EfT@��E�E]��U���E�\E$�E�@�fT�� �E�\E,fT��@�E�\E4fT��@]���������U���Mf(��Y���XU�YM�\��U�E]�����U���M���f(��XU$�E�Y��YM$�\��M�f(��XU,�Y��YM,�\��M�Pf(��XU4�Y��YM4�\��P]��U���E�e]������U���E$�\E�E� �E,�\E�@�E4�\E�@]�������������U���EW�f/��Uvf/�v
�M�E]��^��E�E]�������������U���MW�f/��U4vf/�v(���^��Uf/��],vf/�v(���^��ef/��]$vf/�w(��^ËE� �P�H]�������������U���0�oE����� �~Ef�@�E�P�����oE$����� �~E4f�@�E�P�����UЃ��E����M��Mf��Qf�H����������]������U���0�oE����� �~Ef�@�E�P�)����oE$����� �~E4f�@�E�P�����U���E؋��M��Mf��Qf�H����������]������U���0�oE����� �~Ef�@�E�P�����oE$����� �~E4f�@�E�P�����U���E����M��Mf��Qf�H����������]������U���0�oE����� �~Ef�@�E�P�)����oE$����� �~E4f�@�E�P�����U���E����M��Mf��Qf�H����������]������U���U�E$�XU�XE,�XU�XE4�Yh��Yh�f/�v�E���f� �@]ËEW�f� �@]�������������U���M$�U,�]4�\M�\U�\]����E�X��X��X���P�X]���������U���M$�U,�]4�XM�XU�X]����E�\��\��\���P�X]���������U��E �� H��   HtuHt;�E�M�Y���Y8��X��E�Y��X��M��E���]��oE�~U(�f�f/��E�w�M�f/�vbf(��M��E���]��E�XE�XE�Yh��E��E���]��E�M�YX��Y���X��E�Y��X��M��E���]�����������U����u,�oe���]$��� f�X������M���E�E�]��U��\��\��\��Y��Y��Y��X��X��X�f�� f�X��]��������������U���MW�f/�v��]����f/�r�^@��M�E]��X ��^��(�����U �E�E]��U���MW��@���f/��% ��-���5��v�E��T���f/�r�^��M��;�X��^�(�(��9U �@��% ��-���5���E�W��Mf/�v(��6���f/�r�^��"�X��^�(�(���T �@�f(�W��Uf/��M�w<���f/�r	(��^��%�X �����^��(��T �M��E� �E��H�@��]������U���MW���f/�r�M��E���]�(��x��0T �E��E���]�����U����MW�f/��x��M�s(�(���S �x��E�W��Uf/��U�s(�f(���S �E�W��Mf/�s(��x��S f(ȋE�E��@�E���@��]���U�����MQ�@�@�Ѓ�]��������U������4�@S�]��V�@`Wj �Ћ�   �����   �I V���X� =�   ��   �����V�@�@T�Ћ��Mܡ��Q�u��@�@�С���M܃��@Qj�M̋��   Q���Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M���@Q�M�@x�Ћ������E�P�I�I�ѡ���M�Q�@�@�Ѓ�Fu<�����W�@�@`�Ћ�G�������3�����EP�I�I�у���_^[��]Ëu��������������U���SVW�}����   �]���$    ����ϋ��   �@��;���   =�m u~���x ����tq������� ��uV�E��E�    Ph�  ���E�    ��  ����M�Q���   �@X��SP�k������M������Q���   � uW�Ѓ����W� ����u�����ϋ��   �@4��SP�(�������u*����ϋ��   �@(�Ћ����%���_^3�[��]��Ѓ�_^�   [��]������������U��M��VW�  ����ty�}��$    ����� ��uV�E��E�    Ph�  ���E�    ��� ����M�Q���   �@X��WP�{������M������Q���   � u�Ѓ����g� ����u�_3�^��]��Ѓ��   _^��]����������U��fnE��������} �YEt�E��E��$�s_ �]��,E�����]��E��E��$�4^ �]��,E�����]������U����M�V�q� �E�Phacpihbyek�N� ����M���@j haqpi���   �Ћ��M�#u蔆 ��^��]��������������U���x  ����E�����E��E���   f.�����D{�M����^��   �E��U���   f.�����D{�E����^��   �E��M���   �U�E���E�}���   �M��$�HR �} ��   �M��I �E؋U���   �������E���   �������M��*�������U��*B�������E�P�M�Q�U�R�M�M �*E��*M��^��\������^������E�\��   �YE��M��*E��*M��^��\������^������U�\��   �YE��E�@��	  �M��`Q�UR��X���P��Y  ����X����Y�X�����h����Y�h����X����$�(` ���]��E�f.�����DzH�M������`���f/��v�U����B��E����@�C  ��X����^EЃ��$�}d  ��ݝ�����������^(��M����f/�h���v�U����\�E� �M�U��\��   �E� �M���   f/��v)�U���f/v�E� �X���M��<�U���f/��   v'�E� f/��v�M��\���U��E� �YE��M���`����^EЃ��$�c  ��ݝ�����������^��U�B�E�@�\���M�X��   fWP��YE��U�B�  �E��`P�MQ��p���R�W  ����p����Y�p����M��YM��X����$�
^ ���]��E�f.�����DzH�E���� ��x���f/��v�M����A��U����B�   ��p����^Eȃ��$�_b  ��ݝ8�����8����^(��E� ���f/E�v�M����\�U���x����^Eȃ��$�@b  ��ݝ ����� ����^�����\ȋE�H������Q�����R�E� �Y(����$�\ ������Y������M�YA�X���U�\��   �YE��E� ����Y�����M�YA�X���U�\��   �YE��E�@�  �M��`Q�UR��@���P��U  ����@����Y�@�����P����Y�P����X����$�\ ���]��E�f.�����Dz�M�����  ��@����^E����$�`  ��ݝ�����������^(��U����f/�P���v�E����\ �M��U�E��\��   �M��U���   f/��v)�E���f/ v�M��X���U��<�E���f/��   v'�M�f/��v�U��\���E� �M��YE��U���H����Y���\���E�X��   fWP��YE��M�A��  �U��`R�EP������Q�T  ���������Y���X���U�\��   �YE��E� �������Y���\���M�X��   fWP��YE��U�B�o  �E��`P�MQ�U�R�S  ���E��`P�MQ�U�R�T  ���E��$�_  ��ݝ ����� ������M��$��������^  ��ݝ����������f/�����vj���E��$�^  ��ݝ�������������M��$��0����^  ��ݝ(�����0���f/�(���v	�E�    ��E�   �h���E��$�P^  ��ݝ�����������M��$������%^  ��ݝ���������f/�����v	�E�   ��E�   �E�E�}� t�}���   �}��T  ��  ���f/E�v6�E�fWP��Y���X���M�\��   �YE��U��,�E��Y���X���E�\��   �YE��M��E��Y���\���U�X��   fWP��YE��E�@�J  ���f/E�v/�E��Y���X���M�\��   �YE��U�B�5�E�fWP��Y���X���E�\��   �YE��M�A�E��Y���X���U�\��   �YE��E� �   ���f/E�v.�E��Y���X���M�\��   �YE��U��4�E�fWP��Y���X���E�\��   �YE��M��E��Y���\���U�X��   fWP��YE��E�@�M���   ��t	�   �[�Y�E� f/��r>�M���f/r-�U�Bf/��r�E���f/@r	�E�   ��E�    �E���]ÍI L �M aN /G �M H 1J �����������̡����  � 8���;��@����������U�����M��� �@VW�u�@(Q�Ћ�����}W�I�I�ы��WV�A�@�С���M�Q�@�@�С�����ϋ@�@<�Ћu;���   ������M�Q�@�@�С���M�j j�h|��@Q�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M��� �@�@<�Ћ��j�j�W�Q�M�P�BL�С���M�WQ�@�@�С���M�Q�@�@�С���M�Q�@�@�Ћ�����Q�ϋR<��;��6�����_^��]���������������U������0�@VW�}�@W�С��j j�hx��@W�@��j�E�h�  P�p����ȡ��WQ�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�@�E�jj
P�������M���Q�@�@�С���M�Q�M�Q�@�@�С���M����@�@<�Ћȡ��j��@�@Lj�VQ�M��С���ϋ@�@<�ЋȍU���j�j�R�@Q�ϋ@L�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@��j�E�j
P�,������M���Q�@�@�С���M�Q�M�Q�@�@�С���M���8�@�@<�Ћȡ��j�j�V�@Q�M��@L�С���ϋ@�@<�ЋȍU���j�j�R�@Q�ϋ@L�С���M�Q�@�@�С���H�E�P�I�ы���E�P�I�I�у���_^��]��U������0�@VW�}�@W�С��j j�hx��@W�@��j�E�jP�3����ȡ��WQ�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�@�E�jjP��������M���Q�@�@�С���M�Q�M�Q�@�@�С���M����@�@<�Ћȡ��j��@�@Lj�VQ�M��С���ϋ@�@<�ЋȍU���j�j�R�@Q�ϋ@L�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@��j�E�jWP��������M���Q�@�@�С���M�Q�M�Q�@�@�С���M���8�@�@<�Ћȡ��j�j�V�@Q�M��@L�С���ϋ@�@<�ЋȍU���j�j�R�@Q�ϋ@L�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ��} ��   ����M�Q�@�@�С���M�j j�h���@Q�@�ЍE�P�O������M���Q�@�@�С���M�Q�M�Q�@�@�С���M���$�@�@<�Ћȡ��j�j�V�@Q�M��@L�С���ϋ@�@<�ЋȍU���j�j�R�@Q�ϋ@L�С���M�Q�@�@�С���H�E�P�I�ы���E�P�I�I�у���_^��]�����U�����M����@Q�@�С���M�j j�h���@Q�@�ЍE�P��T ����M�Q�@�@�Ѓ���]���������������U�����M����@Q�@�С���M�j j�h���@Q�@�ЍE�P�T ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h��@Q�@�ЍE�P�AT ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�L�E�P��S ����M�Q�@�@�Ѓ���]��U�����M���`�@VQ�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h ��@Q�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���MЃ�4�@�@<�Ћ��j�j��Q�MQP�MЋBL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�ЍE�j P����������E�P�I�I�ы���A�M�Q�M�Q�@�С���M����@�@<�Ћ��j�j�V�Q�M�P�BL�ЍE�P�uR ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M��@�@Q�С���M�Q�@�@�С���M�j j�h��@Q�@�ЍE�P�K���������E�P�I�I�ы���A�M�Q�M�Q�@�С���MЃ�@�@�@<�Ћ��j�j�V�Q�M�P�BL�ЍE�P�~Q ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ�^��]���U�����M��� �@Q�@�С���M�j j�h ��@Q�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M��� �@�@<�Ћ��j�j��Q�MQP�M��BL�ЍE�P�P ����M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���]����������U���SV3�h�   Sh���]��N h���� h�   h�  h��h�� �@� �� ��tzh��h�   h�j�sC ������t���G �س�3�����M�Q�@�@�С���M�j j�h8��@Q�@��V�E�   h    P�Z{ �� ��t���3���t����E�P�I�I�у���^[��]������������U��� j#h/� �G ������   ����M�Q�@�@�С���M�j j�hȴ�@Q�@�С���M�Q�@�@�С���M�j j�hԴ�@Q�@��hƖ� j �E�P�E�Ph0� h/� ��� ����M���@�@Q�@�С���M�Q�@�@�Ѓ��   ��]���������������U��E���   ����V��i�|  ���b �$�|b �E^�    �@   ��]ËE^�    �@   ��]ËE^�    �@   ��]ËE^�    �@�   ��]ËE^�    �@    ��]ËE^�    �@x   ��]ËE^�    �@   ��]ËE^�    �@
   ��]ËE^�    �@    ��]�(���EЋMfE�P����E��6  �E^��]�(`���p����Mf�p���P����E��R6  �E^��]�(��E��MfE�PW��E��*6  �E^��]�(p���@����Mf�@���P�����P�����5  �E^��]�(���E�MfE�P����E���5  �E^��]�( ��E��MfE�P�(��E��5  �E^��]�(0��E��MfE�P����E��m5  �E^��]�(����X����Mf�X���P� ���h����75  �E^��]�(����(����Mf�(���P�H���8����5  �E^��]ËE^�     �@    ��]��_ ` #` 8` M` b` w` �` �` a �` �` >a ta �a �a �a 1b gb   	
��������������U���\V�$P �����h&� �A�ʋ@T�Ћ�����  �M��+i ����O �����Vh&� �A�ʋ@D�ЍM��di ��O �����h&� �A�ʋ@T�Ћ���u^��]á���M��E�   �E�   Q���   �@8�Ћ�����Q��PhM  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��PhR  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��RhN  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����QP�B4��hO  �С���M�Q���   � �С���M��E�   �E��   Q���   �@8�Ћ�����Q��PhP  �B4�С���M�Q���   � �С���M��E�   �E�    Q���   �@8�Ћ�����Q��PhQ  �B4�С���M�Q���   � �С���M��E�   �E�x   Q���   �@8�Ћ�����Q��PhS  �B4�С���M�Q���   � �С���M��E�   �E�   ���   �@8Q�Ћ������ҋA��Rh]  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��PhT  �B4�С���M�Q���   � �С���M��E�   �E�
   Q���   �@8�Ћ�����Q��PhU  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��Rh\  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��Ph_  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��RhZ  �΋@0�С���M�Q���   � �С���M��E�   �E�    Q���   �@8�Ћ������ҋA��Rh[  �΋@0�С���M�Q���   � �Ѓ�(���E�fE��M����P�E��/  ����M�Q���   �@@�Ћ�����Q��Ph^  �BH�С���M�Q���   � ��(`��E����M�fE����P�E��.  ����M�Q���   �@@�Ћ�����Q��PhW  �BH�С���M�Q���   � ��(��E����M�fE�W�P�E��H.  ����M�Q���   �@@�Ћ�����Q��PhX  �BH�С�����   �M�Q� �С���M��E�   �E�   Q���   �@8�Ѓ��M�fn�������QhY  ��f�E��E��@�@H�С���M�Q���   � ��(p��E����M�fE����P�E��{-  ����M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE����P�E��-  ����M�Q���   �@@�Ћ�����QP�BH��h�  �С���M�Q���   � ��( ��E����M�fE��(�P�E��,  ����M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(0��E����M�fE����P�E��C,  ����M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE�� �P�E���+  ����M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE��H�P�E��s+  ����M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � �Ѓ���^��]����������U�������u0�m(f(��]f(��e�\��}�\��M �\��\��Y��Y��$�Y��X�f(��Y��X�W��^�f/�w.f/��v�]�e �f(��Y$�Y��X��X�(��\��\��Y��Y��X�(��I6 �$�$��]��������������U����j �u�@@�@8�Ѓ�]�������U��M��t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ�]�3�]���������������[c ������    ������������h���Fc �����    �=�� th���5 �����    ���������U���������VW���   �@X�Ћ��u�����   �}��������   �΋@(�Ћ���tK�u���j-��1 ����M�Q�@�@�С���M�j j�h4��@Q�@�С���M�Q�@�@�Ѓ�����M����   �@L�ЍE�P��e ���u����r���_^��]������������̡�����V3����   �@X�Ѕ�t�I ���F���   �ȋR(�҅�u��^�����U�������V���   �@X�Ѕ�t�u;�t������   �ȋB(�Ѕ�u�3�^]ø   ^]�������̡�����S���   �@X�Ћ؅�tzVW�3�W���� ����t;������   ����RX�҅�t ��I ;�t#������   �ȋB(�Ѕ�u�j j W���Y� G��c|�����ˋ��   �@(�Ћ؅�u�_^[��������U��=�� u3�]�VW�u�����������}3��ϋ��   ���   �Ѕ�~M��I �����V���   ���   �Ћ��P���   ����Bh�С����F���   ���   ��;�|������_�   ^]�����������U��=�� tuW�}��tl�����V���   ���   �С��������   �@X�Ћ���t9���$    ����V���   �ϋ��   �С���΋��   �@(�Ћ���u�^_]��������������U������ �@VW���   �@��V�С��j j�h(��@V�@�Ѓ��� 3ɋ�����VD��@�@�С��j j�h,��@V�@�Ѓ�諌 3ɋ�����VD��@�@�С��j j�h0��@V�@�Ѓ��� 3ɋ�����VD��@�@�С��j j�h4��@V�@�Ѓ��_� 3Ʌ�D�hh�h�   h�j��/ ���� ��t����3 �T��3�����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M�j j�h8��@Q�@��V�E�Pj j �E�Ph� �� ����M���@�@Q�@�С���M�Q�@�@�С������@V�@�С��j j�h@��@V�@�Ѓ��� 3ɋ�����VD��@�@�С��j �@�@j�hD�V�Ѓ��>� 3ɋ�����VD��@�@�С��j j�hH��@V�@�Ѓ��(� 3ɋ�����VD��@�@�С��j j�hL��@V�@�Ѓ��� hh�3Ʌ�h�   h�jD��5. ���� ��t���E2 �T��3�����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M�j j�hP��@Q�@��V�E�Pj j �E�Ph� �~ ����M���@�@Q�@�С���M�Q�@�@�С������@V�@�С��j j�hX��@V�@�Ѓ��'� hh�3Ʌ�h�   h�jD��:- ���� ��t���J1 �T��3�����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M�j j�h\��@Q�@��V�E�Pj j �E�Ph� �~ ����M���@�@Q�@�С���M�Q�@�@�С������@V�@�С��j j�hd��@V�@�Ѓ�茄 3ɋ�����VD��@�@�С��j �@�@j�hh�V�Ѓ��֔ 3ɋ�����VD��@�@�С��j j�hl��@V�@�Ѓ��� hh�3Ʌ�h�   h�jD���+ ���� ��t����/ �T��3�����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M�j j�hp��@Q�@��V�E�Pj j �E�Ph� �} ����M���@�@Q�@�С���M�Q�@�@�С������@V�@�С��j j�hx��@V�@�Ѓ��� 3ɋ�����VD��@�@�С��j �@�@j�h|�V�Ѓ��� 3ɋ�����VD��@�@�С��j j�h���@V�@�Ѓ�號 3ɋ�����VD��@�@�С��j j�h���@V�@�Ѓ��3� 3ɋ�����VD��@�@�С��j j�h���@V�@�Ѓ��]� ��3Ʌ�D���_^��]������������VW�9� ������m� ���#�袩 ���#��� ���#�茲 ���#���� ���#��6� ���#�諽 ���#��� ���#��� ���#��J� ���#��� ���#���� ���#��)� ���#��^� ���#���� ���#��� ���#���� ���#��2� ���#���� ���#��\� ���#��� ���#���� ���#��{� ���#��p� ���#��%� ���#��� ���#��O� ���#�脺 ���#���� ���#���� ���#��� ���#��� ���#��� ���#��� ���#���� ���#��l� ���#��a� ��_�#�^���������VW�	� �������� ���#���� ���#���� ���#���� ���#���� ���#���� ���#��� ���#��  ���#�� ��_�#�^�������������U��U��u��+ �Ѕ���   ���h-� R�AL���   �ЋЃ���to���Vj R�A@�@8�Ћ�����tSW�����  ����tDW���&�  ����t6S�]j ���C� ��t�����V���   ���   ��W���� ����u�[_^]�������U������VW���   ���   ���u�E�P�)����u��M�3���9}�   E��>� PWVh+� ��� ���M��ƛ ����M�Q���   ���   �Ѓ�_^��]�������U��E��dt8HtHu+�����t!Pj�s ]��Et�����tj��s �   ]Ë����t����q�@P�@�Ѓ���u�3�]���������Vh��jeh�j�& ������t����r ����F    �5���
���    h�  hR� j h@{ �G4 ���   ^��������������V�5����t �������r V�" �����    hR� j �4 ��^�����U����SV�u�@@�ً@,�Ћ�������Q��j h�  �Rp�ҋ��j h�  �A�΋@4���u����� ^�   []� �U��E��t	�E]��Y ���V�u���   �N�@��-�� t��t��&t�F    3�^]� �F   �   ^]� �����U��W��� t.�O��t'���j Q�@@�@8�Ѓ��ȋj �u�w�RD_]� ���SV�u�@@V�@,�Ћ�����΋؋��   �RT�ҋ��j Ph�  �Q�ˋBl�Ћ���u�G^[3�_]� ����΋��   �@��=�� u�w�   ����΋��   �@��=�� ���u!�@��j h�  ���   ���  P��  �6���   �΋@��=մ u0�����h  h�  �@���   ��P�K�  ����P� � �G�O���H������j Q�@@�@8�Ѓ��ȋj �u�w�RD^[_]� ���������V��N��t���j Q�@@�@8�Ѓ��ȋ�v�RL^� �����U��V��N��t-���j Q�@@�@8�Ѓ��ȋj �u�v�uV�RH��^]� �EW�^ �@]� ���U��Q���VW�}�@@W�M��@,�Ћ���������   �ϋRT�ҋ��j Ph�  �Q�΋Bl�ЋM��j �Z� � -�  tL��t�u�M��u�u�uW�W _^��]� ��tP����΋��   �@��3�=մ _����^��]� ��t&����΋��   �@��3�=�� _����^��]� _3�^��]� �U���E   V��t�U�B    �B    ��u�f� �U�F�B�B   �u���u�u�uR�V ^]� �������������U�����M�@�@ ��=neoa��   VW=ateg��   �% �Ѕ���   ���h-� R�AL���   �ЋЃ���t���j R�A@�@8�Ћ�����te���e�  ����tXW�����  ����tJS�]j ����� ��t�����V���   ���   ��W���B� ����uϋE[_^�    �@   ]ËE_^�    �@    ]ËE�    �@   ]��U���hS�]VWS��| ������E�P�I�I�ы���A�M�QV�@�С���M���@�@<�Ѕ��  ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�SQ�@�@(�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M̃�8�@�@<�Ћ��j�j��Q�M�QP�M̋BL�ЍE�P��+ ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ�3��q  �}W�u{ ������E�P�I�I�ы���A�M�QV�@�С���M܃��@�@<�Ѕ�����@u~�@�M�Q�С���M�j j�h���@Q�@�ЍE�WP�D P�E�P�E�P�t  P�.+ ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ�83��  �u�΋@<�Ѕ���   j VS�ƃ ������   ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E�P�E�P�E�P�E�P�  ��P�E�P�  P�J* ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ� 3��  ����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E��M�P��S j j �0�E��uj PS�mS ���M�������T ����M�Q�@�@�С������ti�@�M�Q�@�С���M�j j�h���@Q�@�ЍE�P�E�P�E�P�  P�C) ����M�Q�@�@�С���M�Q�@�@�Ѓ�,3��  �@���j h�~ ���   �Ћ�����Q�M܋R<�҅���   ���E܋�P�F  �5��������Ѓ���t����A�M�Q���   �M���F ����M�Qj�M��@�@8�С���M�Q���� V�@�M��@8�С���M�Q���V�@�@8�С������P�EP���� P�B4�С������P�E�P���� P�BD�ЍM����F �U����M�Q����@�@8���� V�С���M�Q���V�@�@8�С������P�EP���� P�B4��G���@�����d|0j h��M��@  �E�P�' ����M�Q�@�@�Ѓ�3��������Wh�~ �@�@4�о   ����M�Q�@�@�Ѓ�����E�P�I�I�у���_^[��]����������������U�����M��4�@SQ�@�С���M�j j�h,��@Q�@��j �E�Ph-� �� ���M���Q�Ë@�@�С���M��$�@Q�@�С���M�j j��@�@��t,h<�Q�ЍE�P�& ����M�Q�@�@�Ѓ�3�[��]�hh�Q��j j h�  hд j�E�Ph-� �� ���M���Q�Ë@�@�С���M��4�@Q�@�С���M�j j��@�@��t,hp�Q�ЍE�P��% ����M�Q�@�@�Ѓ�3�[��]�h��Q��j j j hp� j �E�Ph*� �}O ���M���Q�Ë@�@�С���M��4�@Q�@�С���M�j j��@�@��t,h��Q�ЍE�P�l% ����M�Q�@�@�Ѓ�3�[��]�h��Q��j �E�Ph)� �)~ ���M���Q�Ë@�@�Ѓ�$�����������M�Q�@�@�С���M�j j�h���@Q�@�ЍE�Ph@� h�.  h�� �������M���Q�Ë@�@�Ѓ�(���;���j h���M��E  �E�Ph�� h�.  h�� �m������M���Q�Ë@�@�Ѓ��������j h���M���  �E�Ph�� h�.  h�� �%������M���Q�Ë@�@�Ѓ��������j h���M��  �E�Ph�� h�.  h̴ ��������M���Q�Ë@�@�Ѓ����c���j h���M��m  �E�Ph� h�.  h�� �������M���Q�Ë@�@�Ѓ�������j h���M��%  �E�Ph� h�.  h�� �M������M���Q�Ë@�@�Ѓ��������j h ��M���  �E�Ph`� h�.  hʴ �������M���Q�Ë@�@�Ѓ��������j h��M��  �E�PhP� h�.  h�� �������M���Q�Ë@�@�Ѓ����C���j h��M��M  �E�Ph�� h�.  hѴ �u������M���Q�Ë@�@�Ѓ��������j h��M��  �E�Ph � h�.  h�� �-������M���Q�Ë@�@�Ѓ��������j h ��M��  �E�Ph � h�.  h�� ��������M���Q�Ë@�@�Ѓ����k���j h(��M��u  �E�Ph�� h�.  h�� �������M���Q�Ë@�@�Ѓ����#���j h0��M��-  �E�Ph�� h�.  h�� �U������M���Q�Ë@�@�Ѓ��������j h<��M���
  �E�PhP� h�.  h�� �������M���Q�Ë@�@�Ѓ��������j hD��M��
  �E�Ph�� h�.  h�� ��������M���Q�Ë@�@�Ѓ����K���j hP��M��U
  �E�Php� h�.  h�� �}������M���Q�Ë@�@�Ѓ�������j h\��M��
  �E�Ph�� h�.  h�� �5������M���Q�Ë@�@�Ѓ��������j hh��M���	  �E�Ph� h�.  h�� ��������M���Q�Ë@�@�Ѓ����s���j hp��M��}	  �E�Phе h�.  hϴ �������M���Q�Ë@�@�Ѓ����+���j h|��M��5	  �E�PhP� h�.  h�� �]������M���Q�Ë@�@�Ѓ��������j h���M���  �E�Ph� h�.  h�� �������M���Q�Ë@�@�Ѓ��������j h���M��  �E�Ph� h�.  h�� ��������M���Q�Ë@�@�Ѓ����S���j h���M��]  �E�Ph�� h�.  h�� �������M���Q�Ë@�@�Ѓ�������j h���M��  �E�Ph�� h�.  hմ �=������M���Q�Ë@�@�Ѓ��������j h���M���  �E�Ph0� h�.  hT� ��������M���Q�Ë@�@�Ѓ����{���j h���M��  �E�Ph@� h�.  hN� �������M���Q�Ë@�@�Ѓ����3���j h���M��=  �E�Ph � h�.  hִ �e������M���Q�Ë@�@�Ѓ��������j h���M���  �E�Ph � h�.  hO� �������M���Q�Ë@�@�Ѓ��������j h���M��  �E�Ph � h�.  hʹ ��������M���Q�Ë@�@�Ѓ����[���j h���M��e  �E�Ph�� h�.  hش �������M���Q�Ë@�@�Ѓ�������j h���M��  �E�Ph�� h�.  h�� �E������M���Q�Ë@�@�Ѓ��������j h ��M���  �E�PhP� h�.  hU� ��������M���Q�Ë@�@�Ѓ��������j h��M��  �E�Ph�� h�.  h״ �������M���Q�Ë@�@�Ѓ����;���j h��M��E  �E�Ph0� h�.  hQ� �m������M���Q�Ë@�@�Ѓ��������j h ��M���  �E�Ph� h�.  hԴ �%������M���Q�Ë@�@�Ѓ��������j h,��M��  �E�PhP� h�.  hд ��������M���Q�Ë@�@�Ѓ����c���j h4��M��m  �E�Phк h�.  hP� �������M���Q�Ë@�@�Ѓ�������Vh<�h�   h�h�  �� ����t���L  ���3�j h��M���  j h��M���  j ht��M���  �E�P�M��MD V�M�Q�0�E�j Ph&� �V_ ���M������FE ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���tj h���  h<�h�   h�j � ����t���<  ���3�j hX��M��'  j h��M��  j h���M��	  �E�P�M��}C V�M�Q�0�E�j Ph�� �^ ���M������vD ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���tj h����   h<�h�   h�j�J ������t���Z �T��3�j hx��M��Q  j h���M��B  V�E�Pj j �E�Ph� ��] ����M�Q�@�@�С���M�Q�@�@�Ѓ� �M�j h����  hP� �E�Ph+� �T� ���M̡��Q�Ë@�@�Ѓ�j ��t2h���M��  �E�P� ����M�Q�@�@�Ѓ�^3�[��]�h��M��  j h��M��w  j j �E�Ph� j �E�Ph.� �Jx ���M̡��Q�Ë@�@�С���M�Q�@�@�Ѓ�$��u�j h,��M��  j hh��M��  hƖ� h/� �E�P�E�Ph� h'� �]� ���M̡��Q�Ë@�@�С���M�Q�@�@�Ѓ� 3�����^[��]�������U��V�u��V�    �F    ������   �@�Ѓ���^]� ���������������U��V�u��V�    �F    ������   �@$�Ѓ���^]� ���������������U����V��V�@�@�С��V�u�@�@�Ѓ���^]� �U����V��V�@�@�С���uj��@�uV�@�Ѓ���^]� ������������U����   V���Z h\���<���� ��F    �F    �� Phl���t����� Php��M�� P�E�P�r1 ��P�E�P�E ��P��X���P�5 ��P�E�P�( ����X����: �M��2 �M��* �M��" ��t���� ��<���� �=�� u�^I j j��M䣠�Q����E �M��� ��^��]������������V��� �N�,��
   ��^�������U��QSVW���Bh �K���������KD�����Kx�����ˍ��   �G   �C�Kj jh���P8�CD�KDj jh���P8�Cx�Kxj jhp��P8_^��[��]���������VW���wX ����w �`�W�NN�F(O`Op��   ��   ��   ��   ��   Ǉ�      Ǉ�       Ǉ�   ����Ǉ�       Ǉ�       Ǉ�      Ǉ�       Ǉ�   ����Ǉ�       Ǉ�       Ǉ       Ǉ      Ǉ      Ǉ      Ǉ  ����Ǉ  �����  �(  �H����F�>�>����G�ǉw�_^�U���SVW����
 ���s���V�@�@�С���{ W�@�@���5 �C�M���Q�@�@�С���M�j j�hP��@Q�@�С���M�VQ�@�@�С���M�Q�@�@���=5 �C�M���Q�@�@�С���M�j j�h`��@Q�@�С���M�WQ�@�@�С���M���D�@Q�@�Ѓ�_^��[��]��������������V���x� ������F8W�����F@�FH   �FL�F\�Fl�F|���   ���   ǆ�       ^�����V���� (�W��X�����V`Vp��   ��   �F4    FP�F8   W��F<    �F`ǆ�      ( ��FxW�f�Vp���   V@f֎�   f֖�   ^������������VW���� �O�l��d �O�GT��\ ��_^�����̡��V��V���   ���   �Ѓ��    ^���������������V�񍎰   W����`��U j �Nx�Fx ��tY �=�� th����D ���Nx��T j �ND�FD ��EY �=�� th���D ���ND�T j �N�F ��Y �=�� th���D ���N�xT _��^��c ���������������U���   �M�y8�iXf(��A@�YAP�q(�Q �Y��E�f(��M��\�f(��A�YIP�E�(��YQ@�Y��M�(��U��Q0�\��E�(��]��qH�Y��Y���x����M��\��E�(��Y�W��u��e��X�(��Y��X�f.џ��Dza�EW�HH H0H@HP� (���@(���@0f�HW�f�H(f�H@����@Hf�HX��]�����^��q�E�(��Y�(��YA@�if(��	�Y�(��YQP�E�f(��Yq(�\��Yi (��\��\��e��Y}��YA0�Y��X��E��\E��Y��X��E��\E��Y}��Y��}�(��\��\��o�x����Y}��X��oE��\��X��U��\U��o]��Y��Y}�f(��Y��I0�Y��X��Ya@�X��m��Y��Y���x����u��E��E�(��Y��YQX�E��E��Y��E�(��YAX�\�f(��YA(���YY(�Y��\��Y��YIP(ƋE�YA@f��\��E��YA8�Y��\��oE��YA �Y��E�f(�f��YAP�ou��\��u��oE��q0�Yq �Y��E��E��YA8�\��o�x����Y��m��E��oE��M�f�� �oE�f��@�E�f��oE��p �`0f��X@�@P��]���������������U��M�U�;u$�A;Bu�A;Bu�A;Bu�A;Bu3�]ø   ]�������U��M�E�I��`�A0�X�YʋE�Y��X	�X��AH�Y��X��A8�Y���I �Y��XI�X��AP�Y��X��A@�Y��H�I(�Y��XI�X��AX�Y��X��H]����������������U����V�uV�@�@�С��V�u�@�@�С�����΋@�@<�Ћ��j�j��u�Q��P�RL�ҋ�^]������������U��M�E�I�`��A0�X�E�Y��Y��X��AH�Y��X��A8�Y���I �Y��X��AP�Y��X��A@�Y��H�I(�Y��X��AX�Y��X��H]��������������U��V��j � ��MS �=�� th���> �����N �Et	V��� ����^]� ����������U��V���P���� �Et	V�� ����^]� ���������U��V���(��Ϯ �Et	V�s� ����^]� ���������U��V���н蟮 �Et	V�C� ����^]� ���������U��V���u �Et	V�� ����^]� ���������������U��V������?� �Et	V��� ����^]� ���������U��V��N<�4���t�� �F<    ����� �Et	V�� ����^]� ����U��V��� ��ϭ �Et	V�s� ����^]� ���������U��V�����蟭 �Et	V�C� ����^]� ���������U��V���к�o� �Et	V�� ����^]� ���������U��V���@��?� �Et	V��� ����^]� ���������U��V���d��� �Et	V�� ����^]� ���������U��V�����߬ �Et	V�� ����^]� ���������U��V�����诬 �Et	V�S� ����^]� ���������U��V������� �Et	V�#� ����^]� ���������U��V������O� �Et	V��� ����^]� ���������U��V��N�������� �Et	V�� ����^]� �����U��V���U����Et	V�� ����^]� ���������������U��V���`��?K �Et	V�c� ����^]� ���������U��V���H�菫 �Et	V�3� ����^]� ���������U��V���Ŀ�_� �Et	V�� ����^]� ���������U��V��F��P�) �FP�) ����H�F P�A�С���H�FP�A�Ѓ������ �Et	V�� ����^]� U��V������Ϫ �Et	V�s� ����^]� ���������U��V�����蟪 �Et	V�C� ����^]� ���������U��V���x��o� �Et	V�� ����^]� ���������U��V������?� �Et	V��� ����^]� ���������U��V������� �Et	V�� ����^]� ���������U��V���ܷ�ߩ �Et	V�� ����^]� ���������U��V����诩 �Et	V�S� ����^]� ���������U��V������� �Et	V�#� ����^]� ���������U��V������O� �Et	V��� ����^]� ���������U��V���,��� �Et	V��� ����^]� ���������U��V���(��� �Et	V�� ����^]� ���������U��V����迨 �Et	V�c� ����^]� ���������U��V�����菨 �Et	V�3� ����^]� ���������U��V������_� �Et	V�� ����^]� ���������U��V��� ��/� �Et	V��� ����^]� ���������U��V���$���� �Et	V�� ����^]� ���������U��V�����ϧ �Et	V�s� ����^]� ���������U��V��N4����t����@ �@T���F4    ��肧 �Et	V�&� ����^]� ������������U��V���D��O� �Et	V��� ����^]� ���������U��V������ �Et	V��� ����^]� ���������U��V���h���� �Et	V�� ����^]� ���������U��V�����迦 �Et	V�c� ����^]� ���������U��V��N �  ���;� �Et	V�/� ����^]� �����U��VW���O�GT���L �O�2U ���K� �Et	W��� ����_^]� ����U��V��N�T��L ����T �Et	V�� ����^]� ���������������U��V�������A �Et	V�� ����^]� ���������U���Mf/��r��]����f/�r��]�(��� �E�E]���U����E��� �E��E���]�����U����EfT@��E��E���]��U���SVW��� � �Ѕ�t7���h-� R�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3�����M�Q�@�@�С���M�j j�h���@Q�@�ЍE�P� ����t~���j����@V�@�С���M�VQ�@�@�Ѓ����U� �ˋ��H ���+�����P��G ���+�����P��� ��������$�� V���O� �   �3�����E�P�I�I�у���_^[��]���������Vh��h6  h�j@��� ������t%���i� ������P��F4   �F8^�3�^��������Vh��h�  h�j`�y� ������tE���� (����F8�(�����FH   �FL    �FP�FX   �F\   ^�3�^��������Vh|�h�   h�jx�	� ������tY��詢 W��нN8��NHNX�Fh   W��Fl   �F8(�f�NH����FPf�N`�Np^�3�^����Vhp�jbh�jP�� ������t%���,� W����N8��W��F8f�NH^�3�^�����������Vh|�h
  h�j@�9� ������t&���١ �4����F4   �F8    �F<    ^�3�^�������Vh|�h�  h�j<��� ������t��艡 � ����F4    �F8    ^�3�^��������������Vh��h2  h�jP�� ������t5���9� W�����F4    ���F8   �F@�FH   �FL    ^�3�^��������Vh��h�   h�jL�9� ������t;���٠ �к���F4   �F8   �F<   �F@    �FD   �FH   ^�3�^��Vh|�hc  h�j@��� ������t%���y� ������@��F4    �F8^�3�^��������Vh��h�  h�j`�� ������t@���)� ( ���F8�d�W��FP   �FH�FT   �FX   �F\    ^�3�^�������������Vh��h  h�j`�� ������tA��蹟 ������F8W��F@������FH    �FP�FX   ^�3�^������������Vh��h�  h�jH�� ������t,���I� �x�������F8�F@   �FD    ^�3�^�Vh��h�   h�jh�Y� ������t'����� W����F8��(�FHFX^�3�^������Vh��h�  h�jH�	� ������t%��詞 ���������F8�F@    ^�3�^��������Vh��hQ  h�jX�� ������t+���Y� (����F8�H�W��FP   �FH^�3�^��Vh|�hR  h�h�   �f� ������tI���� W��ĿF8���FP    �FHFX�Fx    �Fh����Fp���   ^�3�^�h�h�  h�j0��� ����t������3�����������Vh��h;  h�jH��� ������t%���i� ���������F8�F@   ^�3�^��������Vh|�h�  h�h�   �v� ������tS���� (�W�������F4    �F8   �F<    �F@�NH�FPNX�FhNp��   ^�3�^�������Vh��h�  h�jH��� ������t,��虜 ������x��F8�F@    �FD   ^�3�^�Vh��j`h�jX�� ������t;���L� W�����F@������F4    �F8    �FH�FP   ^�3�^�����Vh|�h�  h�j4�I� ������t���� �����^�3�^������������Vh��hs  h�j4�	� ������t��詛 �ܷ��^�3�^������������Vh|�jh�j@��� ������t%���l� ��������F4    �F8^�3�^�����������h��h�  h�h�   �w� ����t������3��������Vh��hB  h�j4�I� ������t���� �����^�3�^������������Vh��h�  h�jP�	� ������t#��詚 (�����,�F8�FH    ^�3�^����������Vh��jh�j4�� ������t���\� �(���^�3�^���������������h��h  h�h�   �w� ����t�������3��������Vh��h�  h�jX�I� ������tB���� W�����F8������F4    �F@�FH   �FL   �FP    ^�3�^�����������VhX�j.h�j��� ������t����� ������F    �F    ^�3�^�Vh��h(  h�jP�� ������t:���9� ���������F8�F@   �FD   �FH   �FL    ^�3�^���Vh��jh�j@�<� ������t&���ܘ � ����F4    �F8   �F<   ^�3�^����������Vh��h  h�j`��� ������t@��艘 (����F8�$�W��FP   �FH�FT   �FX   �F\    ^�3�^�������������Vh��h%  h�j8�y� ������t���� �����F4    ^�3�^�����Vhp�jh�j8�<� ������t���ܗ �����F4    ^�3�^��������Vh��h�  h�j4��� ������t��虗 �D���^�3�^������������Vh��jh�h�   �� ������t7���Y� W���F8��FH�FX(�F`(P�Fp^�3�^������Vh��jah�j�\� ������t���l� �h���^�3�^���������������Vh,�h�  h�j4�� ������t��蹖 �����^�3�^������������Vh,�jXh�j��� ������t���L� ����^�3�^���������������Vh��jh�j�� ������t���� �H���^�3�^���������������U��VWh��juh�jH���V� ������t:���v �u��PV�� V�O �x��+ W��G@    �G8�G_^]� _3�^]� �����������U�������   ���   ]�����������U���V���t ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���P�yt ����M�Q�@�@�Ѓ���h�� �t ���"u h�� ���t h�� ���t h�� ���t h�� ���t ����t hô ���ot ����t h�� ���\t h�� ���Pt ���t h�� ���=t ���t ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���P�s ����M�Q�@�@�Ѓ���h�� ��s ���Ft hƴ ����s hĴ ���s hŴ ���s ���t hǴ ���s hɴ ���s ����s h�� ���s ���Is ����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E���P��r ����M�Q�@�@��h�.  �5? ����P�r hd� ���s he� ���s h�� ����r ���r h�.  ��> ����P�zr hf� ����r hy� ����r hg� ���r hh� ���r hi� ���r hj� ���r h}� ���r hk� ���zr ���Cr h�.  �y> ����P��q hl� ���Rr hm� ���Fr hn� ���:r ���r h�.  �9> ����P�q ho� ���r hp� ���r hq� ����q hr� ����q hs� ����q h{� ����q ht� ����q hv� ���q ���q h�.  �= ����P�Bq hw� ���q hx� ���q h� ���~q ���Gq h�.  �}= ����P�q h�� ���Vq h�� ���Jq h�� ���>q h�� ���2q hz� ���&q h�� ���q hu� ���q h�� ���q h�� ����p h�� ����p h~� ����p h|� ����p h�� ����p ���p ���p ����M�Q�@�@�С��j j��@�@�M�h�Q�Ѓ��E���P�p ����M�Q�@�@�Ѓ���h&� �_p h'� ���Sp h(� ���Gp h)� ���;p h*� ���/p h+� ���#p h,� ���p h-� ���p h.� ����o h/� ����o ���o ���p ^��]�U���V���Bo ����M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ��E���P�9o ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  �zo ����M�Q�@�@�Ѓ����o ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  �!o ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  ��n ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  �n ����M�Q�@�@�Ѓ����n ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E�P���m ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  ��m ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  �m ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E�Ph�  ���Bm ����M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  ��l ����M�Q�@�@�Ѓ����m ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  �l ����M�Q�@�@�Ѓ����l ����M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E���Ph�  �Al ����M�Q�@�@�Ѓ�����k ���l ^��]�����������U���W���? ��   SV������G�-0 ����D0 �M�_W���Gfn�fn��������G�O ��tI�,�P�,�P�� �M�wVS�8� �M�� ��]��M��Y��O(���Y��^[_��]� ��U��E��wT�$�T� ��  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]Ã��]�� 	� � � � O� %� ,� O� 3� O� :� A� H� ����U��E��wQ�$��� 3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø
   ]Ã��]ÍI �� �� �� �� �� �� �� �� �� �� �� �� �� �� ����U��E��wT�$��� �@  ]øB  ]øC  ]øD  ]øE  ]øF  ]øG  ]øH  ]øI  ]øA  ]øL  ]Ã��]�B� I� P� W� ^� �� e� l� �� s� �� z� �� �� ����U������  �EV��W�t$�    �~P �@    �@�����@    �@    �W  ��� �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��vP���A�  ������NTj h\  �R�|$���   �ҋ���NTjhY  �R�D$d���   �҉D$X����  ��I ���j W�@@�@8�Ѓ����t$;}�y  �|$\ ��   �L$��$�   WP�I �n�  ��$�   ��$�   �Y����P�D$$��$�   �Y���D$<�� �L$��$�   ��$�   � �X�\d$ �\\$8�AH�i(�Y��Y��Y��Y��A8�X�f/���  �X�f/���  �Q0�A@�X�f/���  �X�f/���  ���3��@d�Ѕ��y  �����W�@\�Ѕ��S  �L$W脉 �D$,���=  �t$��$   W�t$�� P����  jc�t$0���o ��$  P�D$|�D$D���  �ЋD$X�T$0�o�D$H���c  �D$p�2   �\D$HW���$�   ��$�   ��$�   fT@��Y����$�   ��$�   ��$�   �,���2��Xl$PLȃ������l$Pfn��������$�   ��$�   ��$�   �D$(�L$(fn��������o�$�   ��$�   ��$�   �X���$�   �(��Xt$`f��X��L$(W��D$���o�t$H� �ă�����$�   f�� �ă���f�� �����$�   P��� �D$ �   ��$�   �D$8��$�   �D$�o�$�   ��$�   �D$H��$�   E�o�$�   D$`���$    �fnƃ�����L$H���^H��D$���o�L$@� �ă��o�$�   �I ��ă����� ��$�   P�!� ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��l$�D$��$�   �f(��D$�D$`��\��T$h�\���\�f(��\�(��Y��Y��Y��X�f(��Y��X�W��^�f/�w)f/��v�l$f(��(��Y��Y��X��X��L$h�D$`�\��\��Y��Y��X���� �0�f/���  �o�$�   F�o�$�   �o�$�   ��$�   ���]����y  ���q  �D$H�}�L$L�\$P�D$0�D$8�T$@�e�u�D$�D$<�|$p�|$0��m���L$8�L$��D$8�\��\$ �\$T�T$H�T$D��D$8�D$ �d$8��\$H�f(��D$ �\��\��|$0�|$p��L$�Y��D$Hf(��l$H�\�f(��Y��Y��X�f(��Y��X�W��^�f/�v�D$�-f/��v�D$0�\$ �(��Y��Y��X��XD$�\��\��Y��Y��X�f(��� �0�f/�wA�t$���G�@d��;�������|$�D$���pP��� ���|$���I����E_^��]� �M�D$�A�D$,�y_�A���   ^��]� ����������U����S�]V�@@WS�@,�Ћ�������Q��j h�  ���   �ҋ�������   �ˋR��=�� ��   ����   �����V�u�@h�  �@l�ЋЅ�tn���jR�AH���  �Ћ�����؋Q��Vh�  ���   ��;�t8�����Sh�  �@�@4�С���MVhȴ ���   �@��_�F^[]� _��^[]� �������������U������   �ES��VW�\$�{P �    �@    �@�����@    �@    �o  �� �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��sP���p�  ������KTj hU  �R�t$���   �ҋKTj h\  fn��������@���   �D$x�Ћ��|$����  ���j V�@@�@8�Ѓ���;u��  ����   �|$��$�   VP�O 螹  ��$�   ��$�   �Y����P�D$4��$�   �Y���D$�� �GH��$�   ��$�   � �X�\d$0�\\$�o(�Y��Y��Y��Y��G8�X�f/���  �X�f/���  �W0�G@�X�f/���  �X�f/���  ���3��Pd����  ���W�P\���x  W����� �D$D���d  �t$jcP��$�   P�N �]�  W�t$�N �o ��$�   P�D$l��$�   �5�  �]�}�u�o�e�T$P�l$P(��D$X��U����T$0��$�   �l$H�l$x�D$�T$ �T$H��l$(�ol$`�L$((��T$H��U�l$l��D$�\����L$(�T$`�oT$0�\$`�f(��D$0�D$�D$ ��l$0�\��\��D$ f(��\��Y�f(��Y��Y��l$0�X�f(��Y��X�W��^�f/�v�l$(�D$ �=f/��v�l$H�D$�%f(��YT$0�Y��XD$((��D$ �X�f(��\��\��Y��Y��X�f(��� �L$pf/���   �L$P�D$X�\�$�   �\L$x�Y��Y��X��� �Y���L$P�\M�D$`�D$X�\E�Y��Y��X��L� �\$pf(��D$`f(��X�f/�v
�\�f/�w@�t$���G�Pd;��h����|$�D$���pP�} ���t$���7����E_^[��]� �M�D$�y_�A�D$@^�A���   [��]� ���������������U���SV��W�FH�E�ǆ�      ǆ�   �����B� �ȅ�t7���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3ۡ��j ���   �@@�@8�Ѓ����~P ��   ���    ��   ����PT����   ����Pd����   ���j �P\����   ���   j �} ����   P�E���P���   �� ��ur�M�f�f.�����DzW����   f^�E�fE����   �΃���� �E�P������}�u"�oE�E����   ���   �   _^[��]�_^3�[��]��������������U���DSW�}3ۉ]�����  ���h-� W�@L���   �ЋЃ�����  ���SR�A@�@8�Ѓ��E����v  V�u��u���w  �����  9]��   ����M�Q�@�@�С���M�j j�hH��@Q�@�С���M�Q�@�@�С���M�j j�h��@Q�@�Ѓ�(�E܋λ   j$P�ʤ P�E�P�E�P������P�E�P������P�f� ���E��t�E ��t����M�Q����@�@�Ѓ���t����M�Q����@�@�Ѓ���t����M�Q����@�@�Ѓ���t����M�Q�@�@�Ѓ��} t^_3�[��]� �M�WV�~+  j j h�� � � j j h,� �� ���   ^_[��]� _3�[��]� �������VW���� �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��wP���`�  ����tj���q� �wP����x ����u�_^���������������U���,�}�  V����   �u�M��O� ���* ���Phdiem�Q�M�B4�С���M�havem�@�@X�Ћ�M�Q���P@�����Phavem�Q�M싂�   �С���M�Q���   � �Ѓ��E��P�* �M���� �   ^��]� �����������������������������������������������U��E��|SVW��=�  ��   tl=�  �l  ����u��j havem�@���   �Ѓ�d�G  �����j j�@���   ��j P��腶  Ph�� �� ���   _^[��]� j h�� �]� ���   _^[��]� F�������  �$��� ��� ����  jj P�������_^�   [��]� �M���� j h@��M��ɻ��j hH��M�躻���E�P�E�Pj j �M��� ���Mԡ��Q�Ë@�@�С���M�Q�@�@�Ѓ���u7j �E�jP�� ���E��t �L� ��tP�u�����  �EP�� ���M��I� _^�   [��]� �� ����  �������  PQ����  _^�   [��]� ��� ��V���������s  �E����  �M���� j h@��M������j hP��M�豺���E�P�E�Pjj �M���� ���M����Q�Ë@�@�С���M�Q�@�@�Ѓ����*����� �E��t&�u��PV��  ��thBF j�E�P�u�l� ���EP�p� ���E    �M��.� _^�   [��]� ��� ��V�#��������r  �؅���  �=�� th���� �����    ��� SPV�ϣ���+  _^�   [��]� �� ��V����������q  �؅��^  �=�� th���� �����    �� SPV�ϣ����  j SV���M���_^�   [��]� �*� P�E�Q����������� ����  �M��5� j h@��M�����j hP��M�������E�P�E�Pjj �M��C� ���M����Q�Ë@�@�С���M�Q�@�@�Ѓ����p������ �E���h�����芄  ����t�]�V�u��S��  ���� ����u�hBF j�E�P�u�� �EP�� ���E    �M��Y� _^�   [��]� �&� ��S�N����������� ����   �=�� th���G� �����    �%� �Σ���ك  ������   V�5����S�@  ���Y� ����u�_�F^[��]� �� P�̌��������o  ����tn���E� P�M��\����E�P��� ����t:�E���P葟 j Vh�� �4� ����M�Q�@�@�Ѓ��   _^[��]� ����M�Q�@�@�Ѓ�_^�   [��]� 0� � �� c�  � �� �� 	� Y� ������������U���VW��� ����躾 ����E�P�I�I�ѡ���M�j j�h��@Q�@�С���M�Q�@�@�Ѓ��σ}cuT�uVj*觾 ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�Ѓ�j�u�u�R�uVj*�S� ����M�Q�@�@�С���M�j j�h ��@Q�@�С���M�Q�@�@�Ѓ�j�u�u����v ���޽ ����M�Q�@�@�С���M�j j�h,��@Q�@�С���M�Q�@�@�Ѓ�_^��]� �������U����oEVj �������(  � �E�P�� �}�ue�M��E�9�  u9�  tm��  ��  9�  t��  cu��cu3���  ^��]� ��cu����  ���@��  ^��]� ǆ      ǆ  ����ǆ      ^��]� ������U���$SV�uW�}��tRV�' �Ѓ����tB���RW�AT�@�Ѓ���t+���v �Ѕ�t������   �ʋ@��=.� ��  �]$��t8���h-� S�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E��E    �M�]q ���W�E�I@�I,��V�E��r h.� �E���t �����ˉu�Vj,�� ����E�P�I�I�ѡ���M�j j�hP��@Q�@�С���M�Q�@�@�Ѓ�����  ���V�@@�@,�Ћ�������Q���uh�  �Rp���u�h �������0����A��Rh�  �@4��Wj(���_� ����M�Q�@�@�С���M�j j�h\��@Q�@�С���M�Q�@�@�С�����ϋ��   j �u����   �С���u�W�@T�@�Ѓ�����t �E�����   ������   �ȋRx�҃��������W�S�@j�u���@����V�С��VW�@�@�ЋM��h�� ��� �����W�@@�@,���oE���������� u ����]����   �ˋ@L��jW�u������M��P�s �����j S���   ���   �С����Sh�  �@�@p�С���u��u��p������M��P�Fp��_^[��]�U���l���SVW�@@�u�@,�Ћ���u�E�I@�I,�ыu$��3��E�}���I W�
 ��S�B$  ������E�Q�M�j S���   �҅��  �E9E��  j �E��E�    PS�M��E�    ��- �MP�k� �M���/ h.� V�M��� ����  ��t8���h-� V�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E���E�    �M��m h.� �E��q ���E��Pj,赸 ����E�P�I�I�ѡ���M�j j�h���@Q�@�С���M�Q�@�@�ЋM��������   �@@Q�@,�Ћ�������Q���uh�  �Rp�ҋ��Sh�  �A�΋@4���u�u$��j(�� ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С�����M���   j �u��   ��j �E��E�    PS�M��E�    �C, �MP��� �M��B. hK  V�M��D� �E�����   ������   �ȋRx�҃��������W�V�@j�u���@����V�С��VW�@�@�ЋM���h�� �� �����W�@@�@,���oE����������q ������   �M��@L��jWS�<  �M��P�o �����j �u����   ���   �С�����u�h�  �@�@p�Ћu$�}����u�M�S�@�@p�С���M�Q���   � �Ѓ�����M�Q���   � �Ѓ�G�}���H�����_^[��]Ë��   �M�Q� �Ѓ�_^[��]��������������U���SV��W�]��ݻ ����t7���h-� W�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3���� �E�������   ���   �ЉE��E����  ���WP�I|�A$�Ѓ�����   �sP���y  �]������   �I j ���j ��t}������u�j ���   � �Ћ���tJWj,���=� ����A�M�Q�@�С���M�j j�hd��@Q�@�С���M�Q�@�@�Ѓ�����M�W���   ���   �ЋE���pP�h �����_�������M����   ���   �Ѕ�tjS�u��\������j�u��@|�@,�Ѓ��J����M�Q�@�@�С���M�j j�h8��@Q�@�ЍE�j P�� ����M�Q�@�@�Ѓ� ����M�Q���   ���   �ЍE��E�    P�4� ��_^[��]� ��������U��Q���V�u�u���   �u�M��v�I�@�С���u�M��u���   �v�I�@�и   ^��]� ��������������U���S�]W���.  ���h-� S�@L���   �ЋЃ����  ���j R�A@�@8�Ћ�������  �U����  ���h-� R�AL���   �ЋЃ�����  ���j R�A@�@8�Ѓ��E�����  V�� �E���u  ���SP�I|�A$�Ѓ����Z  ����u�u��j ���   � �ЋM�jP�E���� V���#v  ������   ���$    ����uj ���   �ϋ ���u�ȉE��l ����E��u����   �H�Rh�ҡ���ϋ��   �@��-�� t��&uy���W�@@�@,�Ѓ���Sh�  �� �Ѕ�tU����uj ���   �ʋ �ЋM��j j V�j� ����u��I@�I,�ы�����ЋA��Vh�  �@p�ЋuV����d �����������j�u�@|�@,�Ѓ��E�   P�� ����^_[��]� �E3�P�� ����^_[��]� _3�[��]� �����U��E=Ҵ u	�E]�Z �E���   ]�+   �����������U��}�� u���  �   ]� ������U���@SVW���ж �u����w� �  ��d� �7  ���� ��   tD��,� �  ���� �  ���� �  �{P �  V��菑 �   _^[��]� �{P ��  ����Mj h1icM�@���   �Ћ�����Mj h2icM�R���   ��j PWh���h������K� �   _^[��]� ��CK�����z  ���� �$��� h���h������ϴ �   _^[��]� ��芽���   _^[��]� ��� �T  �r  ��x� ��   �  ��~� �  ���e� ����M�Q�@�@�С���M�j j�ht��@Q�@�С���M�Q�@�@�Ѓ��E���jP��a  �����o V�����  P���,  ���� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ��   _^[��]� hG  ���  ���0  ��荮 ����j hD�蜦���Q�����E���jP�7a  �����o hx� ����>  P���v
  ���_� ����j hP��N����P�����   _^[��]� h�� ���  ����  ����� ����M�Q�@�@�С���M�j j�h\��@Q�@�С���M�Q�@�@�Ѓ��EЋ�jP�`  �����o h� ����  P����	  ��詭 ����M�Q�@�@�С���M�j j�hh��@Q�@�С���M�Q�@�@�Ѓ��   _^[��]� ��cdpu��   ��   ���C������   ���� �$��� W�Gz��������   ���5]  ����   9CP��   P���� �   _^[��]� ����Mj h1icM�@���   ��P���ܦ �   _^[��]� jW�f���W��y������t%����\  ��t9CPtP�j ��蝦 j ��� _^�   [��]� ��� ?�  � �� ��          ��� �� "� ��           ���U��E�C����(�]  �$�X� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� �ʴ ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� �̴ ]� �ʹ ]� �ϴ ]� �д ]� �Ѵ ]� �Դ ]� �մ ]� �ִ ]� �״ ]� �ش ]� �N� ]� �O� ]� �P� ]� �Q� ]� �T� ]� �U� ]� �S� ]� ���]� �� � � � � (� 1� :� C� L� U� ^� g� p� y� �� �� �� �� �� �� �� �� �� �� �� �� �� �� Q� Q� Q�  � 	� � � $� -� 6� ?� H� ����U���SVW��� ����؍E�P�R�R�ҋ��j j�h��A�M�Q�@�Ѓ��E���P� ����M�Q�@�@�С���M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ��E���j Pj jj?h�  �l5 ����M�Q�@�@�Ѓ���j �6 jjjj���06 jj���5 j j �E�����j?h�  ���L3 �E����   j �E���PV�3 ���>5 ���4 jjj h�  ���E������3 �E���j �E�P�GP�J3 ����M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ��E���j Pj jjj ��* ����M�Q�@�@�Ѓ��E�������jjj h�  �2 �E���j �E�P�GDP��2 ����M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ��E���j Pj jjj �s* ����M�Q�@�@�Ѓ��E�������jjj h�  �2 �E���j �E�P�GxP�B2 ����M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ��E���j Pj jjj ��) ����M�Q�@�@�Ѓ����3 ����P$����P_^��[��]��������������j jxj h�  �@+ �   �����������U���VW���!	 ������E�P�R�R�ҋ��j j�hX��A�M�Q�@�Ѓ��E���P� ����M�Q�@�@�С���M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ��E���j Pj jj?h�  �}2 ����M�Q�@�@�Ѓ���j � 3 jjjj���A3 jj���2 j j j?h�  ���. h�  W�O�� ���_2 ���H���_��^��]�U���$SVW���� ����KTjhZ  �R�E����   �҅���  �uV��� ��������  ��������� ��@V�@tD�С��j j�hp��@V�@�Ћu��E����VP��  ���P���   �ϋB|�ЍM��B�С��j j�h|��@V�@�Ћu��E܃���VP�̗  ���P���   �ϋB|�ЍMܡ��Q�@�@�Ѓ����� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ���j j W�R� Wj,���ؤ ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@��j �e� ����j W�h  �M����^� ����E�P�I�I�ѡ��j j�h���@�@�M�Q�С���M�Q�@�@�Ѓ���j �� ��_^[��]� _^3�[��]� ���������������U���SV��u��Ω �E��Ʃ �Ѕ�t7���h-� R�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3��u�E��P�If  j �vP���m  �oE�����u�� ���j�vP�@����@V�С���M�VQ�@�@�Ѓ����u赮 �M���j �� ����E�P�I�I�у���^[��]� ����������U���<SV��W�]��ݨ ���}��t:���h-� W�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E����3��u�j�Eċ�P�HU  �sP���f  �]����te��I ������   �΋@��=�� u3���V�@@�@,�Ћ�����ЋA��j Wh�  �@l��;���   �E����pP�fU ����u��u��M�j �vP�   ����ˋ��   �@��=G  tu=�� uc����ˋ��   �@x���oEă���������u�@j�vP��@����V�С��VW�@�@�ЋM���hմ �� ���}�l3�_^[��]� ����ˋ��   �@x���oEă���������u�@j�vP��@����V�С��VW�@�@�ЋM���h�� 覬 ���E��t��E�ύ4��E��P�
W fn΃���ɋ���@�X��X���f���[ ���W�@@�@,�Ћ�������}�Q��Sh�  �Rp�ҋ���M�j hS  �B�IT���   �ЋM���E��P�V fn΋����� �\��E��@����\�����   �E��E܋@��=G  ��   =�� ��  ��  ���$    �j �E��E�    PV�M��E�    �� P���K� �M��� ����M�Q���   �@8�Ѓ���t7�u��oEԃ���SV�u� ������E�� �XP��E��E�������j V�@�@0�С���M�Q���   � ��F�����  �L����E_^[��]� 3����$    ��I V�E�    �E�    �������M���E�j PW�� P���p� �M��� ����M�Q���   �@8�Ѓ���td�ƃ�tp��tk��tf����MjW�@�@0���u��oEԃ���V� �B�����PS�u������E�� �XP��E��E������Mj W�@�@0�С���M�Q���   � ��F���������E_^[��]� ����������VW���7� ����t5���h-� V�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3�V�wP����  j ���������_^�   �������������U���SVW����� ���}��t5���h-� W�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��sP�ȉE��a  ����t9j ���4R ���sP��t�6Q �M���j�u�V�   ����Q ����uʋ}�������   ���   ��WP�E��'w���u�M����I Pj Vh+� ��8 ���M��� ����M�Q���   ���   �Ѓ���j �m� _^[��]�������U���S�]V�uWVS�	  ����]S�@@�@,�Ћ�������Q��jh�  �R0�ҋ�����   �M�@��-�� tv��t	��&��   ��tISj(���v� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ������j h�  �@�@p���   �����j Vh�  �@�@l�ЋȉM��tl��tLQj-���� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�ЋM��������   �@L�ЍEP�T ����tISj-��肛 ����M�Q�@�@�С���M�j j�hȶ�@Q�@�С���M�Q�@�@�Ѓ�����M���   �@L�ЍEP�G� ���} tj j hlcrd��� ��_^[��]� ����U���SVW�}�ى]�����  �E��tF��虚 ����M�Q�@�@�С���M�j j�h|��@Q�@�С���M�Q�@�@�Ѓ�W�ˉ}�^  �؅�tW���1N �M���j �uS�����ޅ�u�]��K��t7������   �@X�Ћ���t!;�u���w ����u��jV���΁ ��ujj ��迁 �]��tIWj-���� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ�����M���   �@L�ЍEP��� ����tF��腙 ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ�j j hlcrd�� ��_^[��]� ������������U��E0�����wQ�$�X3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø
   ]Ã��]Ë� 'Q.<CQQJ5U��E������I�  �$��	3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø
   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø    ]ø!   ]ø"   ]ø#   ]ø$   ]ø%   ]ø&   ]ø'   ]ø(   ]ø)   ]ø*   ]ø+   ]ø,   ]ø-   ]ø.   ]ø/   ]ø0   ]ø1   ]ø2   ]ø3   ]ø4   ]ø5   ]ø6   ]ø7   ]ø8   ]ø9   ]ø:   ]ø;   ]ø<   ]ø=   ]ø>   ]ø?   ]ø@   ]øA   ]øB   ]øC   ]øD   ]øE   ]øF   ]øG   ]øH   ]Ã��]�"	>	��v	�	}	��
BIPWz������������L	h	&-^e����		��E	o	4;ls����		�	�	�	�	)	0	7	S	Z	a	����	���������������U��E������Iww����$�l��  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]Ã��]�KY!(/6=DR�
`g  				



		

 		

   ����������U��W�}��tM����IV���   �@X�Ћ���t2S�]��$    ���I ;�ujSj ���IM j ��� G ����u�[^_]� �������������������U���SVW�}�M�����H ���@  j ���9H ���/  j ����G �E����  �]3�V���G ��tY��tIWj*���^� ����M�Q�@�@�С���M�j j�hԶ�@Q�@�С���M�Q�@�@�Ѓ�jj V����K F��c|��M��Ej PW�E    �E�����`� ������   ��    ��tIVj*���Ғ ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�Ѓ�j�u����u�dK �E�M�@P�E�EPW�E�����ء ����u�_^[��]� ���������U���,SV�u�M�W����  ����I���   �@X�Ћ�����  �]���2G ;��]  j ���F ���L  ���G ���=  j ���F ���,  j ���F �E���  3��I V����E ��tY��tIWj*��覑 ����M�Q�@�@�С���M�j j�hԶ�@Q�@�С���M�Q�@�@�Ѓ�jj V���;J F��c|��M��Ej PW�E�    �E����訠 �����~   ��tIVj*��� � ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�Ѓ�j�u���u�I �E��M�@P�E��EPW�E�����&� ����u��uj ����C ���������_^[��]� �U���pVW���P �  ����GH�OTh�   �@hP  �E؋��   �ЋOTj hQ  fn��������@���   �E��ЋOTjhN  fn��������@���   �E��Ћ�����OTjhO  �R���   ���o_(��3��oG8��W�f(�f(��\O0�\�D��E��M��E�\��E��E�]��\��E��E��U��M���E�f.���]�\��   ��U�\��   ��DzW�fE��U��]���^��^��]��U��U��]��oE���   ����  ���   �X����   ���   �X����   ݇�   �E��w �]�݇�   �E��
w fnU��]��o��   ���f(�fT@�f/��]��E��U�w�E��\�f/�w�E��F�E����X�W��^E�f/��E��E��$v苓 ��d� �U����]��E��YE��]�f(��E�fT@�f/�w�E��\�f/�w�E��A�E����X�W��^E�f/��E��E��$v�� ��� �]��E؃��YE苏�   �E�P�E��C �U�W��M��\�\H�X���X���U��E��E��E��M��E��E��]��E��E��E��U��U��]�f.ܟ��Dzf.ԟ��D��   ��� �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��wP���XP  ��3��E���tej ���tA ��t;�E���P�B �M����E����XM��XE؋�f��M���XG �E��wP���? ����u��}�u�������_^��]� U���  V��W�~ ��  �$� �ȅ�t7���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3��E��u���<  �E���Y  ���j �M�����P�]��j �u���IO  (`��M������fE�Q����������E��BhW  Q�N���   �}��ЍM�QhX  �o ������Q�N�������~@���fօ����(�fE�W��E��@���   �Ѓ��o �� ����~@fօ0����E��Y8�f/���E��E��$v�4� ��� �N���]��E��\��jhY  �,��E����@���   �ЋN�E��E�P�E�P�E�Ph�  �}� fnE�E��p�����NP�E�P�E�P�^�h�  ������fnE�����^�������fnE�����^�������� fnE��p�����^��E�fnE�����^��E�fnE�����^��E����d  ��$    ���j W�@@�@8�Ѓ��E�3����W�R\�҅��  �M�W�> �E����  �������W�u�P�w  �jc�u�� �\������H����@��|����\������H����M�P��P�����P����M��Zw  �e���T����]�� �\�����=����U��\���h����@�2   �\������l�����h����W��M���p�����t�����p������L����\��f(���@����\��]��e�fT@��Y���,ȃ�2Lȋ���fn�����E��E��E��E��E��E��E��E��E�fn������8�����8�����x�����<�����|�����@����E���D����E��}�uw�E��X��Y��������E��X��Y���������x����X��Y��������E��X��Y�������f(��Y�������f(��Y��������}�\�E��\�M�f(�f(��\��\��Y5���Y-���X��X��Y��Y���X�����`�����   9E��   9M��   9}u|�N�� ���P�� �Mč������YM܋�j�u�P���L$�M��YM��$�B%  �oE�j ���ă�� �E�f�@���o� ���� �~�0�����  �U ��t	����   9E$��   9M,��   9}(u|�N�� ���P�� �Mč������YM܋�j�u�P���L$�M��YM��$�$  �oE�j ���ă�� �E�f�@���o� ���� �~�0����  j ���: �N����   h�  �� �Mč������YM܋�j�u�P���L$�M��YM��$�$  �N������P�����P�� ���Ph�  �a� �oE�j ���ă�� �E�f�@���o������ ������t������P��� �Mč������YM܋�j�u�P���L$�M��YM��$�{#  �oE�j ���ă�� �E�f�@���o������ �~������u�f�@���o�X�������� �X  �E�G��c������u�M���7 ���}��������_^��]�, �����������U���@W���O����  V��� �O�E���� �M�E�� c ����Oh�   hP  �B�]苀�   �ЋOj hQ  fn��������@�YE苀�   �E��ЋMfn��E����P�YE��E��%b �Oh�  ��H�YU��YM�fWP��U�fWP��M��k� �u��u��OVj j ��� �O�E�W�PfE��E��� �,E�O�u�Pj P�{� �,E��OPVPj �i� �Oh�  �� �E��M��\��E�f/��r4�u��O�,�VPj P�+� �E��M��\�f/���E�sҋu��E��X�fn�����E�f/�r0�u��O�,�Pj P��� �E��XE�fn�����E�f/�s��E��M��\�f/���E�r0���O�,�PVPj �� �E��M��\�f/���E�s��E��X�fnM�����E�f/�r6��I �O�,�PVPj �?� �E��E��XE�fn�����E�f/�sϋOj�5� �O�E�W�h�  PfE��E��� ����M�Q�@�@�С���M�j j�hD��@Q�@���E����X���Oj �,��E��X�P�,�P�E�P�7� ����M�Q�@�@�Ѓ�^_��]� �����������U��V��~ ��   W�� 3�9~u9~t�   h  �h�  ����� �u���u�u�u�S� ����5���@�@�Ѓ�����   �N0�F,h   QP�v(�v$QPj j �5�����?� ��tdh�  ���� �F,��j HPj j �� �F0��HPj j j �� h�  ���O� �N0�F,IQHPQj ���� �F0�N,HIPQj Q���w� _^]� �U���XSV��W�E��� �]�ËM+��u�}P��+�PQ�M�W�=� �M�j�S� �M�h�  ��� S�]���V�uW�F� �{P tv�ۅ �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��H�sP��t#������   �@X�Ѕ�t;�t���] ��u��CP    �CP����   j���� ���+���P��� (��+���P���ă�� �0�f�@��(`������ V���f�@����@�@�С��j j�h���@V�@�Ѓ��K�T  _^[��]� P�K ������A���sP�K�C�O����o��   ���   ���̃���A���o��   ���   �sP��A�K�0����sP�K�  �sP�K�J  �oCp���K�ă�� ���s\�oC`�sP� ��  �o�  �o�   �E��o�   f~��E��~�0  �E��M���tR�}� �Kth�  ��� �(���E�fE�PW��E��� �,E��KP�,E�P�,E�P�,E�P��� _^[��]� ���������S�܃������U�k�l$���  VW���}� ��  �^� �ȅ�t;���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ���4����
ǅ4���    �K��[ �s���@���Pݝh����Ti  ��@����������Y���KP�E���H����Y���E���2 �K� �\E��E��@�������\E�P��p�����Z ����Oj hT  �@���   �Ѓ��E	   fn�����Y�h���f/���E��E��$v螁 ��w� ��h������Y����]�f/���E��E��$v�d� ��=� �E���Y�����]�f/���E��E��$�E�v�(� ��� ��h������Y8���ݝP���f/���E��E��$v�� ��� �s����ݝ`�����1 (����x������f�x���Q����������E��E��Bh^  Q�O���   ��j V�o �������������~@����E؋@@�@8��������O����fWP�U�j�]��E��U��M���X]���X�p����u��]��U���� ��h����� ����E�f��Y��� ����E��Y�������@���fY������Z �K�d/ �� �������������������� �����t[�O����   h�  ��� ������X�����o� ����O�,�f(��X����P�,�P�,����P�,�P�/� �P���ϋă� �}� t(��� � ��W�� f�@��(�f�� ��f��@��  �o� �������������������X���X���\=���\-��( ��O�]���p����m���x����@�f�E��� �����ta��x���P�� �E��XE��o� ����O�,�f(��X�p���P�,�P�,E�P�,�P�� �o� ����]��m���p����}� f(��E�f(�O�X��Y����X���W��X��u�(��\�(��X��u���8���t(���x����0�f�M��(��� ���x���f�E���ta��x���P��� �E��X�8����O�,���X����XE�P�,�P�,E�P�,�X���P�)� ��p����m��]��o� ����,U��,�R����f��E��E��X��f���@����,�(�f��,ȉ�<�����<����,�Q�M��O)E�P��\����w� �������Q���PP�}� �������O�r  �@��������\��������\��\��Y��Y��Y��X��X��X�������f֝����f���������������tN������P�t� �E��XE�O�,���@����XE�P�,�P�u���\������ �������o������,�`���j ���ă���@����XM�(��e��Xe���\�P���f�X��Q���e���� �0�f�@��f����  �K�E�P�8. ����ЋA�ʋ@<�Ћ������E�P�I�I�у�����   �-`������������������\��@��\��e؃�(��\�����0��Y��Y��Y���@����X��X�P����X�f�H���X�f���`����X���f�`�,��E�P��fЋ���?  ����U��,E�j( ��Y�P(P��X�@����,�P���ă�� �@�f�@���f�X��  f֝�����o�������������tN������P�J� �E��XE�O�,���@����XE�P�,�P�u���\����� �������o������,�`���j ���ă���@����XM�(P��e��Xe���\�P���f�X��Q���e���� ���f�@��f���  �K�E�P�, ����ЋA�ʋ@<�Ћ������E�P�I�I�у�����   �o���������������e�(�f(�f��Y�f(ă��Y��Y���@����X�P���f��f�@����`����X���(f�`�,��E�P��fЋ���=	  �U�W��Y��j�,E��X�@���(�P�,�P���ă�� f�@������f�@�K�U��p' ���������IV�I�ы��VW�A�@�Ћ}������  fnE��O���j�XE��,��u��� �K�f* ����  ����Ojh_  �@���   ��@������+��fn�����Y�h����E��E��$�gw �,E����O��p����X��Pݝh����,�P�,� ����u�P��� �,�h������oE�fn�����\��M��,�fn�����Y���E��E��$��v �]��,E؋Kj Qfn�����X�@����,�fn�����E�����@@�E��XE��@8�,��Ѓ���t;�H0��t4�}� �  �   EU�P�,�h���jZjZj j PPVRQ�O�� �?�O������W�Pf������������� �,�h����U��P�
�OPVR�!� �E��Y���XE��XE��,��u�����Oj h]  �@���   �Ѕ���   �K�E�P��' ����M��@�@<�Ѕ���   �,E�Ofn����P��<����,��E�P��\����a� �E��XE�j�,�P�,E�P���ă��}� ��Vt(P�����(������f�@����@�@�С���M�VQ�@�@�Ѓ�����  �E��XE��,��u�����M�Q�@�@�Ѓ��K������P�3& ����������@�@<�Ѕ���   �,E�Ofn����P��<����,��E�P��\����l� �E��XE�j�,�P�,E�P���ă��}� ��Vt(P�����(������f�@����@�@�С��������VQ�@�@�Ѓ�����  �E��XE��,��u�u��u����E�    ��@d�Ѕ���  3ɋQ�΋@\�Ѕ���  �,E�OfnE����P��<����,��E�P��\����� �}� ��u��,  �M�Q���PX(@��O�������`�fօ������tHh�  ������P��� �E��XEȋOj�,���@����XE�P�X��,�P�E�P�� ����M�Q�@�@����@������X�P����K�u��������E��XE��E���! ( ����o��������@P���ă�� �@�f�@��(�� �0�f�@�,�`����E�P��fȋ����  �9  �M�Q���PX(P��O���������fօ������tHh�  ������P�� �E��XEȋOj�,���@����XE�P�X��,�P�E�P�m� ����M�Q�@�@����@���������X�P�������u��@`������Q�E����XE��E����u��K���  ( ����o��������@P���ă�� �@�f�@���o� �~Ff�@�,�`����E�P��fȋ���  �u��E��XE��,��E����E��@d�ЋM�;��%�����΋@T�Ѕ���  �,E�O��p����X��fnM�P����,�P�,�P�,� ���P�� ��4����E�j P�s��z �ȋE������fn��}� �M����t~( �3�(����o� ������U��X�p���P���Xԋă��\�P���� �@�f�@���0�f��f�@�,�`���P������   �o� ���������jc�X�p���Q�@`���\�P����� ����E��X��E���( �3�9M����o� �����Q���̃�����@�f�A�o� �~Bf�@�,�`����E�P��fȋ������  �O�� �OP�� �OPj j �#� ���������Q�@�@�Ѓ�_^��]��[� �U���8fnEW����V�����Y��f/��E��E��$v��n ���m �M�   �U���]��,E�W�;�L��Nfn�����\��\��oE4�X��X��E��~ED�M��U�f�E؅�tL�E�P��� fnM��ɋNf(��XE��,�f(��XE�P�,�P�,E�P�,E�P�R� �M��U��X���X���oE�N�M�fnM�U�����E��~E,(�f�E��\���\���U��M��t;�E�P�D� �E��XE��N�,��E��XE�P�,�P�,E�P�,E�P�� ^��]�D �����������U������tfnE���SVW���L$H�Y��f/���D$P�D$P�$v�`m ��9l �m�   �\$P�,L$P��f(�;�LȉL$Dfn�����\��,�f(��Xŉ|$0fn����f/��7  � ��}�����]׉T$4f(��\��,�f(��XÉ\$(fn����f/���  �4I�]����ˉL$,�I W��Yڋ��D$<   �D$Hf(��YD$8�\$P�D$`�fnȋ���ɻ   �\��Y��L$X�I fn�����\��Y��X��'j fn����f/�w.�}L tf(��\ �f/�w�T$H�X���T$H��T$H�L$XG�\$PKu��D$8�D$`@�L$<�L$,�D$8�X����^8�f.�����D{v�M�D$h�\M4�L$@P�YʋI�XM4�L$l�M$�\M<�Y��XM<�L$t�M,�\MD�Y��XMD�L$|�ƽ �|$0�\$(�D$@WSW�HS�N� ��\$(�|$0�D$DC�]�L$,� ����m�T$4fn����\$(�L$,fn����f(��X�f/��H�����Gf(��Xŉ|$0���T$4fn����f/������_^[��]�H �������U���4S�ى]��{ �*  �Ek �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3�VW�}��W�(  ������   ���E�VP���BQ  �E܍E��Y����P�E��E��Y���E��� �C(�U��M�� �X�\e��\]��k�Y��Y��Y��Y��C�X�f/�w6�X�f/�w,�S�C �X�f/�w�]��X�f/�wWV��������]�W���| �����2���_^[��]� ���������U���  ��3ŉE�V�uW��� �<  ��u��i P�1�������  �����  ���B ��������Pݝ�����B �Oj��� �������������$hH�P�LK ��W�j jjh�  ���ă���� Vf�@����@�@�С��������j j�Q�@V�@�Ѓ����@  ���������������$hT�P��J �O��j �¿ ��W�Pjh�  ���ă���� Vf�@����@�@�С��������j j�Q�@V�@�Ѓ�����  �M�_3�^��J ��]� ��������������U��V��N��t;�E(P�:� �E �XE�N�,��E�XEP�,�P�,EP�,EP訽 ^]�8 ���U��Q�} W����   �M �Ef/�vf(��f(��](�,��Uf/ډE�vf(��f(�f/��,ĉEw(�f/�SV�,�w(ӋOh�  �,�褹 �E�OPSP�u��� �OVS�uS�ռ �OV�u�VS�Ǽ �u�E��OPVP趼 ^[_��]�( �������������U���`�E�e�UV ���h �X(E�W@�E�e��U��m��]�E��� �&  H�;  ��f(��\�fT@�f/���   ���W����D$���oE�� �ă��oE�� �ă��oE�� ���oE�� �E�P�;q �E �   ;���   fn�����Mfnǃ�����ċ�^��D$���oE�� �ă��oE�� �ă��oE�� ���oE�� �E�P��p �,E��NP�,E�P�,E�P�,E�P�I� E�G�ME�;} �t���_^��]� �,ËNP�,�P�,�P�,�P�� _^��]� ������U��V��N��t#h�  �EP腸 �u8�N�E�u4�u0P�p� ����MQ�@�@�Ѓ�^]�4 �������U��S�ًK��teVWh�  �E0P�3� �������uP�EL�K�P�EH�P�EP�� F��~�G��~֋K�Eh�  P��� �uP�K�E�uL�uHP�� _^����MQ�@�@�Ѓ�[]�L �����U��S�ًK��teVWh�  �u0脷 ��������u<�E8�K�P�E4�P�EP肺 F��~�G��~֋K�Eh�  P�e� �u<�K�E�u8�u4P�P� _^����MQ�@�@�Ѓ�[]�8 �����U���SVW���Pd ��ˉE��Rl������   �u�E�j P�u�E�   �u��1�  ���M�P��� P��荍 �M���� ����M�Q���   � �Ѓ���tm�&!�������j hS  �A�ʋ��   �ЋK���E��P�� �u�fn��������\��@�\�����uW�sf��������� jj���� j �lo ��_^[��]� U���SVW���Pc ��ˉE��Rl������   �u�E�j P�u�M��E�   �u���� P��薌 �M���� ����M�Q���   � �Ѓ���tm�/ �������j hS  �A�ʋ��   �ЋK���E��P�� �u�fn��������\��@�\����W�u�sf���ڢ���� jj���� j �un ��_^[��]� ���������j j h�� �2n ���   � �������j j hɴ �n ���   � �������j j h�� ��m ���   � �������j j h�� ��m ���   � �������j j h�� �m ���   � �������j j h�� �m ���   � �������j j hô �rm ���   � �������j j h�� �Rm ���   � �������j j h�� �2m ���   � �������j j h�� �m ���   � �������h'� �&� ���   � �����������j j hǴ ��l ���   � �������j j h�� �l ���   � �������j j h´ �l ���   � �������j j hƴ �rl ���   � �������j j hĴ �Rl ���   � �������j j hŴ �2l ���   � �������j j hl� �l ���   � �������j j ho� ��k ���   � �������j j hf� ��k ���   � �������j j hy� �k ���   � �������j j hg� �k ���   � �������j j h�� �rk ���   � �������j j hm� �Rk ���   � �������j j hh� �2k ���   � �������j j h�� �k ���   � �������j j hp� ��j ���   � �������j j h�� ��j ���   � �������j j hq� �j ���   � �������j j hr� �j ���   � �������j j hs� �rj ���   � �������j j hi� �Rj ���   � �������j j h�� �2j ���   � �������j j hj� �j ���   � �������j j h{� ��i ���   � �������j j hz� ��i ���   � �������j j h�� �i ���   � �������j j h}� �i ���   � �������j j hx� �ri ���   � �������j j hk� �Ri ���   � �������j j ht� �2i ���   � �������j j h�� �i ���   � �������j j hu� ��h ���   � �������j j hw� ��h ���   � �������j j h�� �h ���   � �������j j h�� �h ���   � �������j j h�� �rh ���   � �������j j hn� �Rh ���   � �������j j hd� �2h ���   � �������j j h~� �h ���   � �������j j h|� ��g ���   � �������j j he� ��g ���   � �������j j h�� �g ���   � �������j j hv� �g ���   � �������j j h� �rg ���   � �������j h,  h�  j�j�h&� j���1� � ��������������U���PVW���M��t4���h-� Q�@L���   �Ћȃ���t���j Q�@@�@8�Ѓ��3��H����  ������   �@X�Ћ�����  �d$ ���2 ��u���n2 ����u�_�F^��]� ���b  ���X  j����������"  �w���4 ���  ����M�SQ�@�@�С���M�j j�hH��@Q�@�С���M�Q�@�@�С���M�j j�hL��@Q�@�Ѓ�(�E�j$P�G@P�E�P�Y{  P�E�P�E�P�V����P�E�P�V����P�ua ���MС��Q�Ë@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���[�;  �w����5 _�   ^��]� �w���]3 ���w��t#�?6 j j h,� �1e ���   _^��]� �7 ����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E�j@P�G@P�E�P�z  P�E�P�E�P�qU����P�E�P�dU����P�+` ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���@�@�M�Q�Ѓ�_�   ^��]� ������Vj h,  h�  j�j�h�� j���� ����tj j h�� ��c ����^� ���U���HSVW����W �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3�(0����sPfE�3�(`�fE��/  �]Ћ�����   �E��E��E��E��E��]��E�j ���$ ��tN�E���P�U �M��E�f/�v�M��E��U�f/�v�E�f/M�v�M�f/E�v�E�G�sP���H ����u��M��U��]��e���e��M��U��\��\��Y���Y���X��X��U��E��E��E��M��E��E��E��E��E��~b��� � �M؋˙+���fn�����\��M���� �M����KP�+���fn�������\��oE�f�� �1 j ��赥 _^[��]���������������� �������������U��} t�M��t�j�]� �����̋IV��t0������   �@X�Ћ���t�����y- ��u���>- ����u�3�^Ë�^á��Q���   �@8�Ѓ������������U��U�A��A�B�B*� �B   �A�B�A �B�   �B)� �B   ]� ��������������U������@�@V�uV�@�С��j j�hx��@V�@�ЋE�����g  �$��R����M�Q�@�@�С���M�j j�h���@Q�@�С���M�VQ�@�@�С���M�Q�@�@�Ѓ� ��^��]� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�VQ�@�@�С���M�Q�@�@�Ѓ� ��^��]� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�VQ�@�@�С���M�Q�@�@�Ѓ� ��^��]� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�VQ�@�@�Ћ���E�P�I�I�у� ��^��]� ��%QQ�Q3R������   ���   ���������������U���dV��M��FH�E�W�fE��y �E��E�    Pjhsuom���E�    �-� ���  ����M�j hxvpi�@���   �ЉE��M����j hyvpi�@���   �ЉE��΍E�P�E�P�ܪ �} ufnE��u����fnE������   �oF8�of(�E�fnE�(����f��X��E�fnE��U��M�����f/��X��E��E��E��E��E�vf(��E��X�f/�vf(��E�f/�vf(��M��X�f/�v(��
�E��U��]�Wɋuf.ٟ��Dz�M���x ��^��]� �^��^���M��F�x ��^��]� ��������U������S�]�M��ˋ��   W�@�Ћ}��P��� ��u_[��]� ���VS�@@�@,�Ћ���������   ���   �щE���u3��   ���S���   �ȋ��   �С����j h�  �@���   �ЉE�M��E��E�_  P�E�    �E�    �� �u��E���P�q� �M����� ��t����A3�9M���@0Qj���С����jh�  �@���   �ЉE�M��E��E�Z  P�E�    �E�    諿 �u��E���P��� �M����#� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�V  P�E�    �E�    �7� �u��E���P�� �M����� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�S  P�E�    �E�    �þ �u��E���P�� �M����;� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�a  P�E�    �E�    �O� �u��E���P�� �M����ǿ ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�U  P�E�    �E�    �۽ �u��E���P�-� �M����S� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�W  P�E�    �E�    �g� �u��E���P�� �M����߾ ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�X  P�E�    �E�    �� �u��E���P�E� �M����k� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�Y  P�E�    �E�    �� �u��E���P��� �M������ ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�\  P�E�    �E�    �� �u��E���P�]� �M���能 ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�]  P�E�    �E�    藻 �u��E���P��� �M����� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�R  P�E�    �E�    �#� �u��E���P�u� �M���蛼 ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�^  P�E�    �E�    诺 �u��E���P�� �M����'� ��t����A3�9M���@0Qj���С����j h�  �@���   �ЉE�M��E��E�T  P�E�    �E�    �;� �u��E���P�� �M���賻 ��t����A3�9M���@0Qj���С����j h�  �@���   �Ћ��E�`  �E��E�    P�M��E�    �ȹ �u��E���P�� �M����@� ��t����A3Ʌ����@0Qj���Ћuj ��5V �M���VW�u�E{ ������E�P���   ���   �у���^_[��]� �������������U��Q���V�u�M��@@�@,�ЋM����j 艻 ����  tuItM��t�u�M��u�u�u�u�  ^��]� �����j h�  �@���   ��3Ƀ�^������]� �����j h�  �@���   ����^�@��]� �����j h�  �@���   �Ѕ�t&�����j h�  �@���   �Ѕ�t	3�^��]� �   ^��]� �����������U��Q���V�u�M��@@�@,�ЋM����j 艺 ����  t,��t�u�M��u�u�u�u� ^��]� j h�  �j h�  ����΋@���   ��^��]� ���U��Q���V�u�M��@@�@,�ЋM����j �	� ����  t:��t,��t�u�M��u�u�u�u�~ ^��]� j h�  �j h�  �j h�  ����΋@���   ��^��]� �����U��Q���S�u�M��@@�@,�ЋM����j �y� �8�  t�u�M��u�u�u�u�� [��]� �����j h�  �@���   ��3Ƀ�[������]� ���������U��Q���V�u�M��@@�@,�ЋM����j ��� ����  t!It�u�M��u�u�u�u�u ^��]� �����j h�  �@���   ��^��]� ��������������U��Q���S�u�M��@@�@,�ЋM����j �y� �8�  t�u�M��u�u�u�u�� [��]� �����j h�  �@���   ��3Ƀ�[������]� �������������������������U��Q���V�u�M��@@�@,�ЋM����j �� ����������   �$�a�����j h�  �@���   �Ѓ�tc�����j h�  �@���   �Ѓ�tE�����j h�  �@���   �Ѓ�t'�����j h�  �@���   �Ѓ�t	3�^��]� �   ^��]� �����j h�  �@���   ��3Ƀ�^������]� �����j h�  �@���   �Ѕ�t������j h�  �@���   �Ѓ��'����u�M��u�u�u�u�e ^��]� ���_|`|`�`������������U��Q���S�u�M��@@�@,�ЋM����j �y� �8�  t�u�M��u�u�u�u�� [��]� �����j h�  �@���   ��[��]� ���U��Q���V�u�M��@@�@,�ЋM����j �	� ����  |`���  ~2���  uP�����j h�  �@���   ��3Ƀ�^������]� �����j h�  �@���   ����^��؋�]� �u�M��u�u�u�u�( ^��]� �U���V�q8�E��  V�E��E�    P�.� ��u�V�E�   �    �B    �    ����E�j ���   �E�PR�I�ы���E�P���   �	�у���^��]� ��������������U���V�u�Q� ������E�P�I�I�ы���A�M�QV�@�С���M����@�@<�Ћu�����V�@�@t2�С��V�H�E�P�I�ы���E�P�I�I�у���^��]� �С��j j�h$��HV�I�ы���E�P�I�I�у���^��]� �����������U�����IW�}���   �@X��u��_]� V�Ћ���t�d$ ���y� ;�tj ���l� ����u�^3�_]� ��^_]� �����̋I��u3�á�����   �@X�������̸�� �����������U�����IW�}���   �@\��u��_]� V�Ћ���t�d$ ����� ;�tj ���l� ����u�^3�_]� ��^_]� �����̡��Q���   �@8�Ѓ�������������VW���GA ������v�I@�I,�у���Wh�  ��h _^��U��E�Q,��E�I0��   ]� ����U���@V�4���( ��M����E�fE�P�(��E��-2������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V����(p��M����E�fE�P����E��1������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V�����(���M����E�fE�P����E���0������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V�T���(���M����E�fE�P�H��E��M0������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V����(0��M����E�fE�P����E��/������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V����(���M����E�fE�P� ��E��/������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ����U��E(�� �P��@]� ��������������̸   ����������̸   ����������̸   ����������̸
   ����������̸   ����������̸I   �����������U��U�B���	w�E(� �@]� R�u� �E]� ������������U���u�u� �E]� �����������U��E��u%�E����p���@�H]� P�u�7 �E]� U��E(� �@]� �������U��E��u�E(� �@]� P�u�� �E]� U��E��
}�E(� �@]� P�u� �E]� ���������������U��E��}�E(� �@]� P�u�v �E]� ���������������U��SVW��3��   ��KV�� ��E�F��
~�M��t�G;�~��ct	_^3�[]� _^�   []� ����U��E��x��~��cu	�   ]� 3�]� �������������U��E��cwJ���k�$��k����q�@@�@,�Ћ�����ЋA��j h8  ���   ��]� �   ]� 3�]� ��kYk�k   ����U��E�� tAHt��bt93�]� ����q�@@�@,�Ћ�����ЋA��j h8  ���   ��]� �   ]� �����������U��E��t��ct3�]� �   ]� ��U�����q�@@�@,�ЋЃ��E��
�G  �$�n���j h�  �A�ʋ��   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� �����j h�  �@���   ��]� 3�]� �I �l�l�lm0mMmjm�m�m�m�mU��3�9E��]� �U��3��}c��]� U��SVW�����3��I �KV�� ��E�F��
|�M�G_^[;�~��ct3�]� �   ]� �����������U��E��x��~��cu	�   ]� 3�]� �������������U����V�q�@@�@,�Ћ����E��H�~  �$�|{���j h/  �A�΋��   �Ѕ��U  j h�  �)  �����j h0  �@���   �Ѕ��(  j h�  ��  �����j h  �@���   �Ѕ���  j h�  ��  �����j h  �@���   �Ѕ���  j h�  �  �����j h  �@���   �Ѕ���  j h�  �u  �����j hG  �@���   �Ѕ��t  j h�  �H  �����j hH  �@���   �Ѕ��G  j h�  �  �����j hI  �@���   �Ѕ��  j h�  ��
  �����j h  �@���   �Ѕ���
  j h�  ��
  �����j hK  �@���   �Ѕ���
  j h�  �
  �����j hL  �@���   �Ѕ���
  j h�  �g
  �����j hM  �@���   �Ѕ��f
  j h�  �:
  �����j h  �@���   �Ѕ��9
  j h�  �
  �����j h  �@���   �Ѕ��
  j h�  ��	  �����j h  �@���   �Ѕ���	  j h�  �	  �����j h  �@���   �Ѕ���	  j h�  �	  �����j h  �@���   �Ѕ���	  j h�  �Y	  �����j h  �@���   �Ѕ��X	  j h�  �,	  �����j h%  �@���   �Ѕ��+	  j h�  ��  �����j h&  �@���   �Ѕ���  j h�  ��  �����j h3  �@���   �Ѕ���  j h�  �  �����j h4  �@���   �Ѕ���  j h�  �x  �����j h  �@���   �Ѕ��w  j h�  �K  �����j h  �@���   �Ѕ��J  j h�  �  �����j h  �@���   �Ѕ��  j h�  ��  �����j h  �@���   �Ѕ���  j h�  ��  �����j h'  �@���   �Ѕ���  j h�  �  �����j h(  �@���   �Ѕ���  j h�  �j  �����j h5  �@���   �Ѕ��i  j h�  �=  �����j h6  �@���   �Ѕ��<  j h�  �  �����j h  �@���   �Ѕ��  j h�  ��  �����j h  �@���   �Ѕ���  j h�  �  �����j h  �@���   �Ѕ���  j h�  �  �����j h  �@���   �Ѕ���  j h�  �\  �����j h)  �@���   �Ѕ��[  j h�  �/  �����j h*  �@���   �Ѕ��.  j h�  �  �����j h7  �@���   �Ѕ��  j h�  ��  �����j h8  �@���   �Ѕ���  j h�  �  �����j h  �@���   �Ѕ���  j h�  �{  �����j h  �@���   �Ѕ��z  j h�  �N  �����j h  �@���   �Ѕ��M  j h�  �!  �����j h  �@���   �Ѕ��   j h�  ��  �����j h+  �@���   �Ѕ���  j h�  ��  �����j h,  �@���   �Ѕ���  j h�  �  �����j h9  �@���   �Ѕ���  j h�  �m  �����j h:  �@���   �Ѕ��l  j h�  �@  �����j h  �@���   �Ѕ��?  j h�  �  �����j h   �@���   �Ѕ��  j h�  ��  �����j h!  �@���   �Ѕ���  j h�  �  �����j h"  �@���   �Ѕ���  j h�  �  �����j h-  �@���   �Ѕ���  j h�  �_  �����j h.  �@���   �Ѕ��^  j h�  �2  �����j h;  �@���   �Ѕ��1  j h�  �  �����j h<  �@���   �Ѕ��  j h�  ��  �����j h  �@���   �Ѕ���  j h�  �  �����j hA  �@���   �Ѕ���  j h�  �~  �����j hB  �@���   �Ѕ��}  j h�  �Q  �����j hC  �@���   �Ѕ��P  j h�  �$  �����j h  �@���   �Ѕ��#  j h�  ��  �����j h1  �@���   �Ѕ���  j h�  ��  �����j h#  �@���   �Ѕ���  j h�  �  �����j hD  �@���   �Ѕ���  j h�  �p  �����j hE  �@���   �Ѕ��o  j h�  �C  �����j hF  �@���   �Ѕ��B  j h�  �  �����j h$  �@���   �Ѕ��  j h�  ��   �����j h2  �@���   �Ѕ���   j h�  �   �����j h  �@���   �Ѕ���   j h�  �   �����j h
  �@���   �Ѕ���   j h�  �e�����j hJ  �@���   �Ѕ�thj h�  �?j h=  �j h>  �j h?  �j h@  ����΋@���   �Ѕ�t'j h�  ����΋@���   �Ѕ�t
�   ^]� 3�^]� ���n*oWo�o�o�op8pep�p�p�pqFqsq�q�q�q'rTr�r�r�rs5sbs�s�s�stCtpt�t�t�t$uQu~u�u�uv2v_v�v�v�vw@wmw�w�w�w!xNx{x�x�xy/y\y�y�y�yz=zjz�z�z�z{{&{/{U��� V�u�F���	wu����M�Q�@�@�С���M�j j�hx��@Q�@�ЍF�P�E�P�VJ  �uP�E�PV�%������H�E�P�I�ы���E�P�I�I�у�0��^��]� ��u5����uV�@�@�Ћ��j j�h��IV�I�у���^��]� V�uV�V� ��^��]� �������������U��U��V�u�� t*HtRV�%� ��^]� ���V�@�@��j j�hD�����V�@�@��j j�h<����V�I�I�у���^]� �����U��U��V�u�� t*HtRV�� ��^]� ���V�@�@��j j�h�����V�@�@��j j�hз���V�I�I�у���^]� �����U��EV�u��u0���V�@�@�Ћ��j j�h���IV�I�у���^]� PV�� ��^]� ����U��EV�u��tPV��� ��^]� ���V�@�@�Ћ��j j�h���IV�I�у���^]� ����U��U��V�u�� tFHt*HtRV�� ��^]� ���V�@�@��j j�h��0���V�@�@��j j�h8�����V�@�@��j j�h0����V�I�I�у���^]� ���������U��EV��
�  �$����Mj h���Z���E^]� �Mj h���C���E^]� �Mj h���,���E^]� �Mj h������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h̸�����E^]� �Mj hԸ����E^]� �Mj hܸ����E^]� �Mj h�����E^]� �Mj h��t���E^]� �uPV�� ��^]� �I ������1�H�_�v���������������U��U��V�u�� tFHt*HtRV�� ��^]� ���V�@�@��j j�h��0���V�@�@��j j�hD�����V�@�@��j j�h<����V�I�I�у���^]� ���������U��EV�u��u0���V�@�@�Ћ��j j�hз�IV�I�у���^]� PV��� ��^]� ����U���0V�u��
��   ����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�VQ�@�@(�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���uV�@�@�С���M�VQ�@�@�С����8�΋@�@<�Ћ��j�j��Q�M�QP�΋BL�С���H�E�P�I�ы���E�P�I�I�у���^��]� V�uV��� ��^��]� ��������U���u�u��� �E]� �����������U���0V�u����   ����M�Q�@�@�С���M�j j�h���@Q�@�С���H�FP�E�P�A(�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���uV�@�@�С���M�VQ�@�@�С����8�΋@�@<�Ћ��j�j��Q�M�QP�΋BL�С���H�E�P�I�ы���E��I�IP�у���^��]� V�uV�� ��^��]� �����U��EV�u��tPV�{� ��^]� ���V�@�@�Ћ��j j�hз�IV�I�у���^]� ����U��EV��H��  �$�8��Mj hh��j���E^]� �Mj hx��S���E^]� �Mj h���<���E^]� �Mj h̸�%���E^]� �Mj h������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h�����E^]� �Mj h ��m���E^]� �Mj h4��V���E^]� �Mj hH��?���E^]� �Mj h`��(���E^]� �Mj hp�����E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h �����E^]� �Mj h �����E^]� �Mj h@��p���E^]� �Mj hP��Y���E^]� �Mj hh��B���E^]� �Mj h���+���E^]� �Mj h������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h ������E^]� �Mj h �����E^]� �Mj h0�����E^]� �Mj hH�����E^]� �Mj hh��s���E^]� �Mj h���\���E^]� �Mj h���E���E^]� �Mj h���.���E^]� �Mj h������E^]� �Mj h �� ���E^]� �Mj h������E^]� �Mj h(������E^]� �Mj hH�����E^]� �Mj hh�����E^]� �Mj h������E^]� �Mj h���v���E^]� �Mj h���_���E^]� �Mj h���H���E^]� �Mj h���1���E^]� �Mj h�����E^]� �Mj h(�����E^]� �Mj hH������E^]� �Mj h`������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h���y���E^]� �Mj h���b���E^]� �Mj h���K���E^]� �Mj h��4���E^]� �Mj h �����E^]� �Mj h4�����E^]� �Mj hD������E^]� �Mj hT������E^]� �Mj hh������E^]� �Mj h|�����E^]� �Mj h������E^]� �Mj h���|���E^]� �Mj h���e���E^]� �Mj h���N���E^]� �Mj h���7���E^]� �Mj h �� ���E^]� �Mj h��	���E^]� �Mj h ������E^]� �uPV�� ��^]� �����ń܄�
�!�8�O�f�}�����م����5�L�c�z�������ֆ���2�I�`�w�������Ӈ���/�F�]�t�������Ј����,�C�Z�q�������͉����)�@�W�n�������ʊ��������U���(���SV���E�    �@Wj�N���   h_  �u���@����+ȡ���j �M��@�NhS  ���   �Ћ��3ۋNShT  �R�E싒�   ��S�u�E	   �E����@@�@8�Ћ�����3���Rd��~���W�P\��tC���G�Pd;�|��u����PT���   E١���M�j h]  �@�I���   �Ћu��t,�E��E�   P����� ����ЋA�ʋ@<���E���u�E� �E�t����M�Q�@�@�Ѓ��}� �   �   ��E��E�P��� ����ЋA�ʋ@<�Ћ�����E�P�Q�R�҃���tG�M� � ��t�U����3�fnE��M�E���_^���[� fn�����@��]� U���X���SV���E�    �@Wj�K���   h_  �]��Ћu@����+ȍE��V�M��P������E��E��Y����P�E��E��Y���E��f� �Kj hT  � �\E��E��@����\EЋ@�Eȋ��   ��3��E�    SVfnȡ����ɋ@@�Y���@8�X8�f(��M��Y���E�f(��X���E��Ћ����EW��� ��� ��t�E��fn�����XE��E����M�j h]  �@�I���   �Ѕ�t,�E��E�   P����� ����ЋA�ʋ@<���E��u�]�E�t����M�Q�@�@�Ѓ�8]t�E��XE��E�E���P�� ����ЋA�ʋ@<�Ћ�����E�P�I�I�у���t�E��XE��E���3��Pd��~*��I ���V�P\���E�t@�E�;u��D؋F�Pd;�|ۃ}c�E�u>�XE��E_^[�\���\E�� �E��XE��XE��\���@��]� �X���M�C��M��XM�_�XE�^[�fn�������YE��X��XE��A��]� ����������̡��jQ�@�@H�Ѓ�������������̡��j Q�@�@H�Ѓ��������������U��E�  ��   ]� ����������̸,�����������̸   @� ��������U��UVW����t4���h-� R�@L���   �Ћȃ���t���j Q�@@�@8�Ѓ��3��H��t.������   �@X�Ћ���t����� ��u���� ����u�3��G���u_3�^]� ��t�P����� ��_�%���?   @^]� ����̸�������������U���VW��� �M���G: �E�P�u�N��g ����M�j Wheert�@�@l�ЍM���v: _��^��]� ������������U���`�MSVW�_� �]����S�@�@�С���MSQ�@�@�Ѓ��E   ����   ���    ����΋��   �@x�Ћ�����E�P�I�I�ы���A�M�QW�@�С���MЃ��@S�@x�Ѕ����tG���   �΋@(�Ћ��MС��Q�@�@�Ѓ���u�����EP�I�I�у���_^[��]� �@�M�Q�@�С���M�j j�h���@Q�@�С���M��uQ�@�@(�Ћ�����E�P�I�I�ы���A�M�QW�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�MQ�@�@�С���M���8�@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�С���M�Q�@�@�M�Q�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�SQ�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M��EQ�@�@�Ѓ��������������̡��Q���   �@@�Ѓ�������������U�����u�u�@�uQ���   �Ѓ�]� ������������U�������@SVW�}�񋀠   ��j hacpi�Ѓ~P �؉^Xj uj h�� �0 ���   _^[��]� ������E    �E�    hxvpi�@���   �ЉE�ϡ��j hyvpi�@���   �ЉE��΍E�P�EP�h fnM��fnE����j �������f���E�P�@O  �����j haqpi�@���   �Ѓ�Ku�M��u�M��t��t��� ��b� j �{ ���   _^[��]� ����������U����SVW�@�ًMj hacpi���   �Ћ�����Mj haqpi�R���   �ҋȋ�у�������cOt�ǽ����   �����$������   ����   ����   QQh�� � ���   _^[]� ��xmtD��dt,��vui��te��ua��u]QQh�� �u ���   _^[]� ���? _^�   []� ��t+��u'��u#QQh�� �; ���   _^[]� ���  t	_^3�[]� j j h�� � ���   _^[]� ���z�S����� ��U������0�@S�]V���   ��Wj hacpi���Ѓ~P ���~Xu&���%  h���h������ �G�_^[��]� hTCAb�M��E�    �E�    �=4 �M��4 ����] ���Phdiem�Q�MЋB4�С���M�j havem�@�@4�С����j hxvpi�@���   �ЉE��ˡ��j hyvpi�@���   �ЉE��΍E�P�E�P�)e �����j haqpi�@���   �Ћ؃�tt��to��tj��d�  ����Mj havpi�@���   ��fnM���fnE���Q�ˋЃ���Q���S���΋����Rf���J  j ���
\ �  �M��fnM�fnE�QP�Ë΃���P���S�������Wf���|<  j ����[ �E��P�vXhsuom�@] ���^  ���    ����M�j hxvpi�@���   �ЉE��M���j hyvpi�@���   �ЉE��΍E�P�E�P��c ����M�j haqpi�@���   �Ћ����j havpi�Q�M䋒�   ��fnM���fnE�����ɋ����f�tg��P�ǃ���PW�����vX���C  j ����Z ����M�jhrdem�@�@4�ЍEЋ�P�X[ �E��P�vXhsuom�5\ ��������Q��P�ǃ���PW�����vX��,F  j ���sZ �FX    �MС��j hrdem�@�@4�ЍEЋ�P��Z j � ���M��1 �M��1 _^�   [��]� ��U���V�uV�� ���V�@@�@,�Ћ�������Q��jh�  �R4�ҋ��������A���$h�  �@,�С����jh9  �@�@4�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M����@Qh<  �΋@8�С���M�Q�@�@�Ѓ��   ^��]� �����U��V�uV�3� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ��������΋@�$h�  �@,�С����jh�  �@�@0�С����j h�  �@�@4�С��������΋@�$h�  �@,�С����jh�  �@�@4�и   ^]� ������������U���V�uV�P� ���V�@@�@,�Ћ�������Q��jh�  �R0�ҡ���M�W�fE�Q�E��΋@h�  �@H�С����jh�  �@�@0��(��M���fE�Q������E��@h�  �@H�С��������΋@�$h�  �@,�и   ^��]� ����������U���u�u� ����u�@@�@,�Ћ�����ЋA��jh>  �@0�и   ]� U���   V�uV�-� ���V�@@�@,�Ћ�������Q��jh�  �R4�ҋ��j h�  �A�΋@4���W� �E��u3���   ����M����W��E��E�W��E�Q(����U��E�    �U��E�    f�M��M��E�f�U��U�豉 �M�E�P襉 ����M��u�E�    �E�    ���   h!D Q�@\�С���M����@Qh�  �΋��   �С���M�Q���   � �Ѓ��   �EP虍 ����^��]� �������������U���V�uV��� ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ��j h�  �A�΋@4�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M����@Qh<  �΋@8�С���M�Q�@�@�Ѓ��   ^��]� ���������U���V�uV�� ���V�@@�@,�Ћ�������Q��jh�  �R4�ҋ����W��A���$h�  �@,�С����jh�  �@�@0���[� �E��tmj���[� �E��t]���P�E�    �E��E�    ���   h�e P�A\�С���M����@Qh�  �΋��   �С���M�Q���   � �Ѓ��EP�� ���   ^��]� ���������������U��V�uV�� ���V�@@�@,�Ћ�������Q��jh�  �R0�ҋ��jh�  �A�΋@0�С����jh�  �@�@0�С����j h�  �@�@4�С����jh�  �@�@4�С����jh�  �@�@4�и   ^]� U���V�uV�P� ���V�@@�@,�Ѓ����� �E��tmj���� �E��t]���P�E�    �E��E�    ���   h�e P�A\�С���M����@Qh�  �΋��   �С���M�Q���   � �Ѓ����������΋@�$h�  �@,�ЍEP�w� ���   ^��]� ��������U��V�uV�s� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ��������΋@�$h�  �@,�С����jh�  �@�@0�С����jh�  �@�@0�С����jh�  �@�@4�и   ^]� U��V�uV�ý ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ����W��΋@�$h�  �@,�С����j h�  �@�@4�С��������΋@�$h�  �@,�С����jh�  �@�@4�и   ^]� �������U��V�uV�� ���V�@@�@,�Ћ�������Q��h�  h�  �R0�ҋ��jh�  �A�΋@4�и   ^]� �����U��V�uV裼 ���V�@@�@,�Ћ��W�Q���$h�  �Q�΋R,�ҡ����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�и   ^]� ������������U��V�uV裻 ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ����j h�  �@�@4�и   ^]� U��V�uV�C� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ��������΋@�$h�  �@,�С����W��΋@�$h�  �@,�С����jh�  �@�@0�и   ^]� �������������U��V�uV蓺 ���V�@@�@,�Ћ��W�Q���$h�  �Q�΋R,�ҡ����W��΋@�$h�  �@,�С����W��΋@�$h�  �@,�С����j h�  �@�@0�С����W��΋@�$h�  �@,�С����W��΋@�$h�  �@,�С����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С���@��j h�  �@0�С��������΋@�$h�  �@,�и   ^]� ������������U����W�u�����   �O�@l�С���u�O���   �@l�и   _]� ����U��V�uV�� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ����jh�  �@�@0�и   ^]� U��V�uV蓸 ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ��jh�  �A�΋@0�С����j h�  �@�@0�С����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С����W��@�@,���$h�  �С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�и   ^]� ���������U��V�uV�ö ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ����j h�  �@�@4�С����jh�  �@�@4�и   ^]� ����������U���V�uV�@� ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ��j h�  �A�΋@0�С����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С���M�Q�@�@�С���M�j j�hT��@Q�@�С���M����@Qh<  �΋@8�С���M�Q�@�@�Ѓ��   ^��]� ��U��]�'� �������U��V�uV�� ���V�@@�@,�Ћ�������Q��jh�  �R0�ҋ��j h�  �A�΋@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����jh�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����jh>  �@�@0�и   ^]� ������������U���V�uV�г ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ��������A���$h�  �@,�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M����@Qh<  �΋@8�С���M�Q�@�@�Ѓ��   ^��]� �����������U��V�uWV�� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ����W��ϋ@�$h�  �@,�С����jh�  �@�@0��3����    �����j �P��M  P�B4��F��|�����jhY  �@�@4��_�   ^]� �U��V�uV�C� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ��������΋@�$h�  �@,�С����j h�  �@�@4�и   ^]� ������������U���V�uV谱 ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ��jh�  �A�΋@0�С����j h�  �@�@0�С����W��΋@�$h�  �@,�С����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С���M�W�fE�Q�E��΋@h�  �@H��( �fE����M��X��E�Q�@��h�  �@H�С���M�W�fE�Q�E��΋@h�  �@H�С����jh�  �@�@0�и   ^��]� ������U���V�uV� � ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ����W��A���$h�  �@,�С��������΋@�$h�  �@,�С����jh�  �@�@0�С����jh�  �@�@4���1} �E��tmj���1 �E��t]���P�E�    �E��E�    ���   h�e P�A\�С���M����@Qh�  �΋��   �С���M�Q���   � �Ѓ��EP��| ���   ^��]� �����U��V�uV�� ���V�@@�@,�Ћ�������Q�$�Q��h�  �R,�ҡ����jh�  �@�@0�С����jh�  �@�@4�и   ^]� ����������U��V�uV�c� ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ��jh�  �A�΋@4�С����jh�  �@�@4�и   ^]� ��U��V�uV�� ���V�@@�@,�Ћ�����0�Q�$�Q��h�  �R,�ҡ��������΋@�$h�  �@,�С����W��΋@�$h�  �@,�С����jh�  �@�@0�С����jh�  �@�@0�С����jh�  �@�@4�и   ^]� �U���V�uV� � ���V�@@�@,�Ћ�������Q��j h�  �R4�ҋ���A�M�Q�@�С���M�j j�hp��@Q�@�С���M����@Qh<  �΋@8�С���M�Q�@�@�Ѓ��   ^��]� ���������������U��V�uV�s� ���V�@@�@,�Ћ�������Q��j h�  �R0�ҋ��j h�  �A�΋@0�С����W��΋@�$h�  �@,�С����W��΋@�$h�  �@,�С����W��΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С��������΋@�$h�  �@,�С���@������@,���$h�  �и   ^]� �����������U��V�uV�#� ���V�@@�@,�Ћ�������Q��j h�  �R0�ҋ��jh�  �A�΋@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����jh�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h�  �@�@0�С����j h/  �@�@0�С����j h0  �@�@0�С����jh  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j hG  �@�@0�С��j hH  �@�@0���С����j hI  �@�@0�С����j h  �@�@0�С����j hK  �@�@0�С����j hL  �@�@0�С����j hM  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С���@��j h%  �@0�С����j h&  �@�@0�С����j h3  �@�@0�С����j h4  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h'  �@�@0�С����j h(  �@�@0�С����j h5  �@�@0�С����j h6  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h)  �@�@0�С����j h*  �@�@0�С����j h7  �@�@0�С����j h8  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С����j h  �@�@0�С���@�@0��j h  �С����j h+  �@�@0�С����j h,  �@�@0�С����j h9  �@�@0�С����j h:  �@�@0�С����j h  �@�@0�С����j h   �@�@0�С����j h!  �@�@0�С����j h"  �@�@0�С����j h-  �@�@0�С����j h.  �@�@0�С����j h;  �@�@0�С����j h<  �@�@0�С����jh  �@�@0�С����j hA  �@�@0�С����j hB  �@�@0�С����j hC  �@�@0�С����j h  �@�@0�С����j h1  �@�@0�С����j h#  �@�@0�С����j hD  �@�@0�С����j hE  �@�@0�С����j hF  �@�@0�С��j �@�@0��h$  �С����j h2  �@�@0�С����j h  �@�@0�С����j h
  �@�@0�С����j hJ  �@�@0�С����j h=  �@�@0�С����j h>  �@�@0�С����j h?  �@�@0�С����j h@  �@�@0�С����jh>  �@�@0�и   ^]� ��������������U���0V��E��MP�oF(ǆ�      ���   �E��oF8�E�臗 �oM�W��o ǆ�      ǆ�       ���   ǆ�       f(�ǆ�   �����\U��\��M�\��E�\�f����   ^��]� ��������̸   � ���������A    �   �A    �������������V���F\    ǆ�       �FX    �����vP�N �FT�����   ^�������������A8���$�^�  �   ���������U���V���B ��u^��]ÍM��� ����M�htxt heman�@�@4�ЍE�Pj�N�	: h�  ����E �M�� �   ^��]������������U���8V��~P ��   �FHW��oN(�E�M�E��oF8P��  �E؉�  �E�f(�  �\V0�\���  QP�N ǆ      �U��E�������@�YM�ǆ      �YE��XM��XE�f��oE��  ��(  ^��]� �������������U��E�A �EH��wb�$�X��A$    �=�A$   �4�A$    �+�A$0   �"�A$@   ��A$P   ��A$`   ��A$p   �A0   �A,   �A(    �E�A   �A]� �I ����������(���������U���0���S�]V�@��Wj hvdpi���   ���Ћ����j hacpi�Q�ˋ��   �҉E��E�    �E    ��suom�S  hTCAb�M���
 �M��
 ���t4 ���Phdiem�Q�M�B4�С���M�j havem�@�@4�Ѓ}���  �����j hxvpi�@���   �ЉE��ˡ��j hyvpi�@���   �ЉE�΍EP�E�P�; j ���F   �3 �F ��t�u�u�jV�v�Ѓ��EЋ�Pjhsuom�{4 ����   �I ����M�j havpi�@���   �Ѕ���   ����M�j hxvpi�@���   �ЉE��MС��j hyvpi�@���   �ЉE�΍EP�E�P�; j ���l2 �F ��t�u�u�jV�v�Ѓ�����M�jhrdem�@�@4�ЍE��P��2 �EЋ�Pjhsuom�3 ���8�������M�j hrdem�@�@4�ЍE��P�2 j ���F    ��1 �F ��t�u�u�jV�v�Ѓ��u����u��P,��t2�~ t3�9F���Fj ���1 �F ��t�u�u�jV�v�Ѓ��M��� �M��� _^�   [��]� _^3�[��]� ��U����V�uW�@��j hvdpi�΋��   ��=byekuV���.���_^]� =suomu6�����j hbdpi�@���   �Ћ�V��t�����_^]� �a���_^]� _3�^]� ���U��Q���E��xP u3���]� S�]��u	3�[��]� W�}��j�k� ��t
_3�[��]� Vj��胘 ���j W�@@�@8�Ѓ��E3����V�R\��t.V���7� ��t"V���+� ;�t!V���� �M�PS�e�����uF��c}�E�^_�   [��]� ^_3�[��]� �������������V��  �t?��   t6�F����  c��u��  ��  �����^���  ��  �����^�3�^��U��� SVW���� �Ѕ�t8���h-� R�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E���E�    �����14 ��3���~V���q4 F;�|��, �E�3��E��E�    �H����   ������   �@X�Ћ���t|��$    �M�� ���!� ���Pheman�Q�M��B8�С���M�Wheert�@�@p�ЍE���PV�83 ���� ��t�M�V��( �u��誶 �M���F�� ��u��u�����3 ���1 j �u���^4 �E�P��+ ��_^[��]������������U�����M����@VW�u�@(Q�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]����U��QSW���G    �L� �؅���   ���h-� S�JL���   �ыЃ�����   ���Vj R�A@�@8�Ћ������~   ���(����E���tpP��艛������tb�I � uHVS���q����t+����΋��   �@�С����j h�� ���   �@���u����� ����u�j j h,� �d� ��^_[��]�����������U���DSVW�}����  ���h-� W�@L���   �ЋЃ�����  ���j R�A@�@8�Ћ؃��]����  �u����  ���h-� V�AL���   �ЋЃ����u  ���j R�A@�@8�Ѓ��E����V  �� �E����-  ���WP�I|�A$�Ѓ����  ���� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�ЋK�����5  ������   �@X�Ћ؅��  �d$ ������u�j ���   � �ЋM�jP�E��\ �u��j,�0� ����A�M�Q�@�С���M�j j�h���@Q�@�С���M�Q�@�@�ЋM��S�W���������  ������u�j ���   � ���u�ȉE��ڏ ����E��u����   �H�Rh���u��Mj,�� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С�����΋��   �@��-�� t	��&��   ���V�@@�@,�Ѓ���Wh�  � �Ѕ���   ����u�j ���   �ʋ �ЋM��j j W�T� �MWj,��� ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���u��@@�@,�Ћ�����ЋA��Wh�  �@p�Ћ}S��臇 ������������Ʊ �u�؅���������j�u��@|�@,�Ѓ����� ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@��j �� j j h�� �� ��(�E��   P�� ����_^[��]� �E�3�P�� ����_^[��]� _^3�[��]� ���������U�������@SVW�}��@ ���Ћ]=fnic�  �~X ��   �~P �t  �����j j�@���   �ЉE�ϡ��j j�@���   �ЉE�΍EP�EP�`1 fnM��fnE���j �������f���E�P�4  ���   P�E�P�d�������t�oE�E��j ���   ���   �( �}� u�E��t	����  �����hfnic�@�@$�С����jj�@�@4��SW����% _^[��]� ����ϋ@�@ ��='  �g  �����j j�@���   �Ѕ��I  �E��ΉE�EP�E�PW�01 �}��   �  �M���  ���j�hG  ���   ���   �Ѕ�u%����Mj�h�� ���   ���   �Ѕ���   j���,1 �����j j�@���   �Ѕ���   �M�����3��E��E    ���~   �����W���   �M���   �Ћ���؋��   �ˋR��=G  t������   �ˋ@��=�� u�~P u��������t�u��S��-���Ej ���j& G;}�|��   _^[��]� j���]0 SW���T$ _^[��]� �����������U����}S��u=�M�E�Pj �E��  �E�    �E�    �H ����C ��tj h&� �� ���u���u�u�� [��]� �������������U���SVW�}�ك���   ��Ҵ ��  ��� ������u�I@�I,�у��E�V��h�  ���p� ����  ��  �I �����j W�@���   �Ћ3PW�6������P�Vp�u�G���  ~��B  �� �ȉE��i� ����E�P�I�I�ѡ���M�j j�hh��@Q�@�С���M�Q�@�@�С���u�@@�@,�ЋM�����u��	j ��F �8��0�����w*�����j W�@���   �Ћ3PW��5������P�Vp�u����  uL�u���W�n� ��t=��  ��I �����j W�@���   �Ћ3PW�5������P�Vp�u�G���  ~͋M��� ����M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�Ѓ��u���u�u�� _^[��]� �������������U��Q�}���E���   ���V�u�@@�@,�Ћ��W�Q���$h�  �Q�΋��   �������W��\$�$h�  V�; ���������΋@�D$W��$h�  ���   ��������$h�  V�� �E���^�u���u�u�?� ��]� ���������U��E��S�]V��W����   =Ҵ �L  �&� �����S�I@�I,�у��؋ˉ]�Wh�  �� ���  ��  �I �����j W�@���   �Ћ��PW�RpG���  ~ٻ  �d$ S�7����������Q�M�j W���   �ҋ��PW�RpC��M  ~��  �� �ȉE��h� ����E�P�I�I�ѡ���M�j j�h��@Q�@�С���M�Q�@�@�С��S�@@�@,�Ћ؃��E�]�j ���C �8�}���0�����w �����j W�@���   �Ћ��PW�Rp�8��������Iw-W�6����������Q��j W���   �ҋ��PW�Rp�}����  u}�u���W�>� ��tn��  ��I �����j W�@���   �Ћ��PW�RpG���  ~ٻ  �d$ S�:6����������Q�M�j W���   �ҋ��PW�RpC��M  ~̋M��4� ����M�Q�@�@�С���M�j j�h ��@Q�@�С���M�Q�@�@�Ѓ��E�]�u��PS賎 _^[��]� ����������U�������@V�uW�@ ������=TCAb��   �����j hdiem�@���   ��=�  ��   �����j hghcv�@���   �Ѕ�u=���������΋@�$havem���   ���]��E�f.�����D{>�����W��΋@�$havem���   �Ѓ����]��E��G8�$��  �u��V��h _^��]� ����������U��]�G, �������U���<  SVW���P ��  �� �ȅ�t7���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3��oEj ���ϋ�� �E�P�  j�wP���-5���oE�E���   H��  Ht#H�f  9E$�]  j��� ��_^[��]�$ �}$ tAj��������P�{��j ���o ������P���   �~{���o ���   _^[��]�$ �} ��  �}  ��  �E�H����  �$�d��M�����  jj j��� �M��� j h���M��d�������M�Qh�� �M�@�@8�С���M�Q�@�@�Ѓ��M�j h���(�������M�Qh�� �M�@�@8�С���M�Q�@�@�Ѓ���D���j h�����������D���Qh�� �M�@�@8�С����D���Q�@�@�Ѓ���T���j h��褿�������T���Qh�� �M�@�@8�С����T���Q�@�@�Ѓ���$���j hx��_���P��t������������t���Qj �M�@���   �С����t���Q���   � �С����$���Q�@�@�Ѓ��M�j h�����������M�Qhô �M�@�@8�С���M�Q�@�@�Ѓ���4���j hx�輾��P�M��C�������M�Qj �M�@���   �С���M�Q���   � �С����4���Q�@�@�Ѓ���d���j h���^�������@��d���Qhɴ �M�@8�С����d���Q�@�@�ЋG�M�j j
Qh���h����p��h ����~j j P��� ���M���� _^[��]�$ �u����+  j �wP����1��jj j���H j �/j j�j �+�u�����  j �wP���1��jj j��� �u��u�Vh���h�������  _^[��]�$ �}$ �Z����} �E���   H��   HtQH��  �u�����  �}�c��  j �E$�E$����PV����  �؅���  �u$��jj V�~ VS��  �u����D  j �wP����0��jj j���a~ V���	�  �(  �}  t;HtUH�  �u����  P���qy ��jj ����   j �~ _^[��]�$ H����  �$�t�j �wP���f0��E�G\   E��oE��G`�Gp_^[��]�$ �}� tmj�2� ��������   ���   �Ћu���j �E$��x ��tj �u$�������	�M$V�����j �u$��h�   �u(�]# �M$����_^[��]�$ �u����  j ���x ��uP�wP���/��jj ��j�,} �oE���ϋ�V� �����_^[��]�$ �}� ��  �u�����  �E�E$�����  �OP�!� �]��M�f.�����DzW�fE��E��E��E��E���E�^��E��E�^��EԋOP�����P�R� �E̋��X �E��@�������XE�P�E���x �E̋M��\ �E��E��\@������P�E��x �]��U��M��\P�\�E��Y��Y��Y��Y��X��X�f/�v�u��c   �E$��E��t=��cu8j�@� ������jcV�oE���ϋ�� � ���_^[��]�$ �]�u���]$j�� ����tX��ct�S���av �E$��tjj S����z jc�u$�S랋M������j@P�z P�=� ��������Q�@�@�Ѓ�_^[��]�$ �L��$�T�����������,�����U���(V��VP����  �M��HtH�  H�~  �}$ ��  �FH�E�P���E�臟 �]�\��   �F`�U�\��   fWP��\�fWP��F`�Fh�\��Fh�Fp�\��Fp�Fx�\��Fx��  �\���  ��   �\���   ��(  �\���(  ��0  �\���0  �E�f.�����D��   W�fE��U��]���   �}$ �u  j �E��P��r���E����\��   �$��=���]��M���fWP�f.�����D�)  �o��   �����vP� ���$�@o �]��E��N �Y���XFH�$��  �oE����   �oE���   ^��]�  �^��^��M؃��E��XˋNP�X�f���^� �oE���   ^��]�  ��u}�~\ t'�oEj ���Fp�ܣ  �oE���   ^��]�  ���    t)�oE���΋�� �.���oE���   ^��]�  ��    t�oE���΋�� �H���oE���   ^��]�  ����U���SV��W�~P ��  �� �؅�t7���h-� S�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3��EHtGHt$H��  9E$��  PPhƴ �� ����  �} ��  j j hǴ ��� ���  �~\ t	j��諢  ��    t(��   t��  ����  ��  ��  ��������   �V  ��覽 ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ������   j*蘽 ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ћ��   ��j���   j �$v ���   ��j*�5� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ����   j���   ���   �u ��趼 ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ�j�vP���F\    ǆ�       ǆ       ǆ�      �6(��j�/� ������   ���   ��j P�E�!����u�M����C0 Pj Vh+� ��W ���M���2 ����MQ���   ���   �Ѓ�_^[��]�  �������U����} VW��tL�}  �
   �NP�   E��E�P�� ����} fn����}�M��\��M��\�XE��E��P�}$ th�}  �
   �NP�   E��E�P衙 ����} fn����}�M��\��M��
�XE��E��oE��NP����� ��� _^��]�  �E��yj j hŴ �~j j hĴ �� ��_�FX    �F\    ǆ�       ǆ       ǆ�      ^��]�  ������������̸   �����������U����   ���V��W�@j �FH�NT���   �E��oF(hT  �u���H����oF8��X����Ћ��+� �ȅ�t7���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3�WɍGf(��}�\�H����vP�   �G    �E��E�f(��\�P���fn�����G�����G    �G    �E��YM��E�f(��M�fWP��E�f(��Y���E��}�����u؅��n  E�E�d$ ���j V�@@�@8�ЋM����E��x���VP�I �w�����x���������Y����P�E��E��Y���E���n �E���x����U�� �\e��X�\]��m�M�Y��Y��Y��Xe��X]��Y��E�� ����E�f/��u��e��]���$����k  (��X�f/���8����R  �� ���f/��@  �X�f/���(����*  �M���h���VP�I �o�����h�����X����Y����P��@�����p����Y����0�����m �M���h�����p���� �X�\�@����\�0����AH�i(�Y��Y��Y��Y��A8�X�f/���   �X�f/�wv�Q0�A@�X�f/�wb�X�f/�wX�M�m�]��E�e�f/��E��e�r,��8���f/�v�U��M�f/�r��(���f/�wU�E����pP��j ���E؅�������?�N  �E�W��M�U�\M��\U�f.ß��D�u  W��  �E��}��X��XM�f(��   �w�e��X��M��]��M��M��E��E��U���E�X��f(��M�X���E�f/�r5�E��X�f/�v&�M�f/�r�X�f/�v�G   ��_^��]� �E܋�P�-n ����ЋA�ʋ@<�Ћ������E�P�I�I�у�����   �E��XE��e��E��E��U��E��E��]��M���E�X��U���M�X��]�E��E�f/��E�r4�E��X�f/�v%�M�f/�r�X�f/�v�   ��_^��]� �M��@T�Ѕ���   �M���X���jc�u�P�I �!����e�� �YE��H�YM��XE��XM��E��U��E���E�X��U��M��]��M���M�X��]�E��E�f/��E�r;�E��X�f/�v,�M�f/�r!�X�f/�v�   ���Gc   _^��]� �M3���@d�Ѕ��J����MV��@\�Ѕ���   �M���X���V�u�P�I �/����e�� �YE��H�YM��XE��XM��E��U��E���E�X��U��M��]��M���M�X��]�E��E�f/��E�r$�M��X�f/�v�E�f/�r
�X�f/�w�MF��@d��;��&����k����   �ǉw_^��]� �^��^��M��U�fE܋u���j ����� ��T���P�����o �@��G�?ui�U�W��E�M�\E��\M�f.ӟ��DzW���^��^��E��M�fE�j ���΋�� ��T���P�e����o �@��G��_^��]� �������������U����   SV��W�u��Z� ���}���t:���h-� W�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E����3ۉ]��=� �E������   ���   �ЉE��E����  ���WP�I|�A$�Ѓ�����  �u��F����C���M��E�������   ���   �Ѕ���  ��舱 ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ���j �vP�M�����W��NTj hR  �@fE����   �Ћ���؋NTj hZ  �R�]����   �҉E����Y  ���3�(0��M�fE싀�   (`�fE����   ���U����   �E��E��E��E��E��U��Eȡ���M�V���   ���   �ЍM�Q���f �M��E�f/�v�M��E��U�f/�v�E�f/M�v�M�f/E�v�EС��F�M����   ���   ��;�|��E��M��U��]���]��E��M��\u��\��Y���Y���X��X��E��M��E��E��E��E��E��E��E��E����3ۋM��]̋��   ���   �Ѕ��  �I ����M�S���   ���   �Ћ؋�Sj(药 �����8���P�I�I�ѡ����8���j j�h���@Q�@�С����8���Q�@�@�С�����ˋ��   �@L�С���M�S���   �@h��Sj,���� �����X���Q�@�@�С����X���j j�h���@Q�@�С����X���Q�@�@�Ѓ����vP��h jj j���h �E��P�d �E���u&�M���E���\M��\E�f����   ��uv�NP��(���P蹍 �NP� �Y���E��@������Y��P�E��g� �U��]��M��@�\U��X�XE��\M��X��X�f��B��uMj��x�����P�}`���E��\E��M��\M���x����X��E��X�fЃ�������ph �vP���6b ���������IV�I�ы��VW�A�@�ЋM��E���P��  �}���Sj(�d� �����H���Q�@�@�С����H���j j�h ��@Q�@�С����H���Q�@�@�Ѓ��E���P�Qf ���S�@@�@,�Ћ�����EԋQ��jh�  �R0�҃}� �  ����ˋ��   �@��-�� t	��&��   ����ˋ��   �@��=�� uhG  �"����ˋ��   �@��=մ ��   h�� �S� ��������   j j V���ʗ Vj,���P� �����h���Q�@�@�С����h���j j�h��@Q�@�С����h���Q�@�@�С�����Mԋ@Vh�  �@p�С����j hҴ ���   �@�С���M�Q�@�@�С�����]̋M�C�]̋��   ���   �Ћu�;���������j�u�@|�@,�ЋM��W�_������X� ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�Ѓ��J����M�Q�@�@�С���M�j j�h���@Q�@�ЍE�j P�Q� ����M�Q�@�@�Ѓ� ����M�Q���   ���   �ЍE��E�    P��� ��_^[��]�������������U��E��
wQ�$���3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø   ]Ã��]ÍI ����������������������U��E��
wT�$�t���  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]Ã��]�"�)�0�7�>�E�L�S�Z�a�h�U��E��H�  �$����/  ]ø0  ]ø  ]ø  ]ø  ]øG  ]øH  ]øI  ]ø  ]øK  ]øL  ]øM  ]ø  ]ø  ]ø  ]ø  ]ø  ]ø  ]ø%  ]ø&  ]ø3  ]ø4  ]ø  ]ø  ]ø  ]ø  ]ø'  ]ø(  ]ø5  ]ø6  ]ø  ]ø  ]ø  ]ø  ]ø)  ]ø*  ]ø7  ]ø8  ]ø  ]ø  ]ø  ]ø  ]ø+  ]ø,  ]ø9  ]ø:  ]ø  ]ø   ]ø!  ]ø"  ]ø-  ]ø.  ]ø;  ]ø<  ]ø  ]øA  ]øB  ]øC  ]ø  ]ø1  ]ø#  ]øD  ]øE  ]øF  ]ø$  ]ø2  ]ø  ]ø
  ]øJ  ]ø=  ]ø>  ]ø?  ]ø@  ]Ã��]Ë������������������������
����&�-�4�;�B�I�P�W�^�e�l�s�z�������������������������������������������"�)�0�7�>�E�L�S�Z�a�h�o�v�}���������������U��W��j�u�O�� �Oj�u� � �   _]� ������U���TVWh+  � ������E�P�I�I�ы���A�M�QV�@��hh�jxh�j脧 ���� ��t��蔫 �l��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M���� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh	+  �� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j�q� ���� ��t��聩 ����3�����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Phɴ �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M���� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���TVWh�*  ��� ������E�P�I�I�ы���A�M�QV�@��hh�jh�j�d� ���� ��t���t� ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M���� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh�*  ��� ������E�P�I�I�ы���A�M�QV�@��hh�jh�j�T� ���� ��t���d� �D��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh�*  ��� ������E�P�I�I�ы���A�M�QV�@��hh�j0h�j�D� ���� ��t���T� ���3�����M�Q�@�@�С���M�j j�h<��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�u� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh�*  �� ������E�P�I�I�ы���A�M�QV�@��hh�jHh�j�4� ���� ��t���D� ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�e� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh+  �� ������E�P�I�I�ы���A�M�QV�@��hh�jTh�j�$� ���� ��t���4� ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�U� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Phô �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh +  �� ������E�P�I�I�ы���A�M�QV�@��hh�j`h�j�� ���� ��t���$� ����3�����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�E� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��v� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh�*  �� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j�� ���� ��t���� ����3�����M�Q�@�@�С���M�j j�h ��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�2� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��c� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���TVWh�*  �~� ������E�P�I�I�ы���A�M�QV�@��hh�j$h�j��� ���� ��t���� ����3�����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�%� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��V� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh+  �n� ������E�P�I�I�ы���A�M�QV�@��hh�jlh�j�� ���� ��t����� �4��3�����M�Q�@�@�С���M�j j�hX��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �w� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��F� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh+  �^� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j�ѐ ���� ��t���� ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�PhǴ �d� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��3� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���TVWh�*  �N� ������E�P�I�I�ы���A�M�QV�@��hh�j<h�j�Ď ���� ��t���Ԓ �L��3�����M�Q�@�@�С���M�j j�hp��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P��� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �W� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��&� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]��������U���TVWh+  �>� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j豌 ���� ��t����� ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P��� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph´ �D� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���TVWh+  �.� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j衊 ���� ��t��豎 ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P��� �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�Phƴ �4� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���TVWh+  �� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j葈 ���� ��t��行 ���3�����M�Q�@�@�С���M�j j�h8��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P�¾ �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�PhĴ �$� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���TVWh+  �� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j聆 ���� ��t��葊 �H��3�����M�Q�@�@�С���M�j j�hl��@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ�(�E��M�P貼 �M�Q�0����@�@�С���M�Q�M�Q�@�@�С���M܃��@�@<�Ћ��j�j��Q�MQP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�Ѓ�����M�@�@<�Ћ��j�j��Q�M�QP�M�BL��W�E�PVj �E�PhŴ �� ������E�P�I�I�ы���A�M�Q�@�Ѓ� �M��� ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���MQ�@�@�Ѓ���_^��]�����U���dVh�� ��� ������E�P�I�I�ы���A�M�QV�@��hh�hR  h�j�r� ���� ��t��肈 �p��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��ҹ V�M�Q�0�E�h   Phl� ��� ���M����˺ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�hs  h�j�2� ���� ��t���B� ���3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h@��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒷 V�M�Q�0�E�h   Pho� �� ���M���苸 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�h  h�j�� ���� ��t���� ���3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h@��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R� V�M�Q�0�E�h   Phf� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh̴ �?� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�} ���� ��t��� �h��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phy� �� ���M����� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� ��� ������E�P�I�I�ы���A�M�QV�@��hh�h  h�j�r{ ���� ��t��� �T��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��Ұ V�M�Q�0�E�h   Phg� ��� ���M����˱ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhT� �� ������E�P�I�I�ы���A�M�QV�@��hh�h{  h�j�2y ���� ��t���B} ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒮 V�M�Q�0�E�h   Ph�� �� ���M���苯 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�h]  h�j��v ���� ��t���{ ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R� V�M�Q�0�E�h   Phm� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �?� ������E�P�I�I�ы���A�M�QV�@��hh�h&  h�j�t ���� ��t����x ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phh� �� ���M����� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhN� ��� ������E�P�I�I�ы���A�M�QV�@��hh�hO  h�j�rr ���� ��t���v ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��ҧ V�M�Q�0�E�h   Ph�� ��� ���M����˨ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�h~  h�j�2p ���� ��t���Bt �T��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�hx��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒥 V�M�Q�0�E�h   Php� �� ���M���苦 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhִ �� ������E�P�I�I�ы���A�M�QV�@��hh�h.  h�j��m ���� ��t���r ���3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h(��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R� V�M�Q�0�E�h   Ph�� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �?� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�k ���� ��t����o ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phq� �� ���M����� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� ��� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�ri ���� ��t���m ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��Ҟ V�M�Q�0�E�h   Phr� �ع ���M����˟ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�2g ���� ��t���Bk ���3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h0��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒜 V�M�Q�0�E�h   Phs� 蘷 ���M���苝 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhʴ �� ������E�P�I�I�ы���A�M�QV�@��hh�h1  h�j��d ���� ��t���i ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R� V�M�Q�0�E�h   Phi� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhO� �?� ������E�P�I�I�ы���A�M�QV�@��hh�hZ  h�j�b ���� ��t����f ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Ph�� �� ���M����� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� ��� ������E�P�I�I�ы���A�M�QV�@��hh�h<  h�j�r` ���� ��t���d � ��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h$��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��ҕ V�M�Q�0�E�h   Phj� �ذ ���M����˖ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhϴ 迺 ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�2^ ���� ��t���Bb ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h ��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒓 V�M�Q�0�E�h   Ph{� 蘮 ���M���苔 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhʹ �� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j��[ ���� ��t���` ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R� V�M�Q�0�E�h   Phz� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhS� �?� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�Y ���� ��t����] ���3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h8��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Ph�� �� ���M����� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhѴ ��� ������E�P�I�I�ы���A�M�QV�@��hh�h  h�j�rW ���� ��t���[ �P��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�ht��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��Ҍ V�M�Q�0�E�h   Ph}� �ا ���M����ˍ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� 迱 ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�2U ���� ��t���BY �,��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�hP��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒊 V�M�Q�0�E�h   Phx� 蘥 ���M���苋 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�hG  h�j��R ���� ��t���W �8��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h\��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R� V�M�Q�0�E�h   Phk� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �?� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�P ���� ��t����T �D��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�hh��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Pht� �� ���M����� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhش ��� ������E�P�I�I�ы���A�M�QV�@��hh�hD  h�j�rN ���� ��t���R �|��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��҃ V�M�Q�0�E�h   Ph�� �؞ ���M����˄ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� 迨 ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�2L ���� ��t���BP �|��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M�蒁 V�M�Q�0�E�h   Phu� 蘜 ���M���苂 ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j��I ���� ��t���N ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��R V�M�Q�0�E�h   Phw� �X� ���M����K� ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhU� �?� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�G ���� ��t����K ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��} V�M�Q�0�E�h   Ph�� �� ���M����~ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh״ ��� ������E�P�I�I�ы���A�M�QV�@��hh�h9  h�j�rE ���� ��t���I �@��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�hd��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M���z V�M�Q�0�E�h   Ph�� �ؕ ���M�����{ ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhQ� 迟 ������E�P�I�I�ы���A�M�QV�@��hh�hp  h�j�2C ���� ��t���BG �d��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��x V�M�Q�0�E�h   Ph�� 蘓 ���M����y ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�hh  h�j��@ ���� ��t���E ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��Rv V�M�Q�0�E�h   Phn� �X� ���M����Kw ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �?� ������E�P�I�I�ы���A�M�QV�@��hh�h�   h�j�> ���� ��t����B ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��t V�M�Q�0�E�h   Phd� �� ���M����u ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhԴ ��� ������E�P�I�I�ы���A�M�QV�@��hh�h  h�j�r< ���� ��t���@ ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M���q V�M�Q�0�E�h   Ph~� �، ���M�����r ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhд 迖 ������E�P�I�I�ы���A�M�QV�@��hh�h  h�j�2: ���� ��t���B> ���3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h<��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��o V�M�Q�0�E�h   Ph|� 蘊 ���M����p ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� �� ������E�P�I�I�ы���A�M�QV�@��hh�h  h�j��7 ���� ��t���< ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��Rm V�M�Q�0�E�h   Phe� �X� ���M����Kn ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhP� �?� ������E�P�I�I�ы���A�M�QV�@��hh�he  h�j�5 ���� ��t����9 �,��3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�hP��@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��k V�M�Q�0�E�h   Ph�� �� ���M����l ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVh�� ��� ������E�P�I�I�ы���A�M�QV�@��hh�h�  h�j�r3 ���� ��t���7 ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M���h V�M�Q�0�E�h   Phv� �؃ ���M�����i ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U���dVhմ 迍 ������E�P�I�I�ы���A�M�QV�@��hh�h#  h�j�21 ���� ��t���B5 ����3�����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M܃�@�@Q�M�Q�@�С���M܃��@�@<�Ћ��j�j��Q�M�QP�M܋BL�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�ЍE�P�M��f V�M�Q�0�E�h   Ph� 蘁 ���M����g ����E�P�I�I�ѡ���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���^��]�����������U�����M��$�@VQ�@�С���M�j j�h���@Q�@��h��j:h�j��. ����$��t���3 ����F    �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�Pe V�M�Q�0��h   Ph&� �W� ���M����Jf ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�hP��@Q�@��h��jEh�j��- ����$��t���2 �,��F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�Pd V�M�Q�0��h   Ph'� �W ���M����Je ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�h���@Q�@��h��jPh�j��, ����$��t���1 �h��F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�Pc V�M�Q�0��h   Ph(� �W~ ���M����Jd ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�h���@Q�@��h��j[h�j��+ ����$��t���0 ����F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�Pb V�M�Q�0��h   Ph)� �W} ���M����Jc ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�h��@Q�@��h��jfh�j��* ����$��t���/ ����F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�Pa V�M�Q�0��h   Ph*� �W| ���M����Jb ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�h@��@Q�@��h��jqh�j��) ����$��t���. ���F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�P` V�M�Q�0��h   Ph+� �W{ ���M����Ja ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�h|��@Q�@��h��j|h�j��( ����$��t���- �X��F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�P_ V�M�Q�0��h   Ph,� �Wz ���M����J` ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]��������������U�����M��$�@VQ�@�С���M�j j�h���@Q�@��h��h�   h�j��' ����$��t���, ����F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�M^ V�M�Q�0��h   Ph-� �Ty ���M����G_ ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]�����������U�����M��$�@VQ�@�С���M�j j�h���@Q�@��h��h�   h�j��& ����$��t���+ ����F   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�M] V�M�Q�0��h   Ph.� �Tx ���M����G^ ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]�����������U�����M��$�@VQ�@�С���M�j j�h0��@Q�@��h��h�   h�j��% ����$��t���* ���F	   �3�����M�Q�@�@�С���M�j j�h��@Q�@�Ѓ��E܍M�P�M\ V�M�Q�0��h   Ph/� �Tw ���M����G] ����E�P�I�I�ѡ���M�Q�@�@�Ѓ���^��]�����������U���(S��W�]��N) �Ѕ�t5���h-� R�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��H��u3��}��������   �@X�Ћ��E�3��E��E���u ���E�P���} ����   V��3��1} ��~Q�( �M؋��NO �E؋�PV��| ���j Wheert�A�M؋@l�ЍM؋��O �E�;�to��F��| ;�|�����M�Q�@�@�С���M�j j�h���@Q�@�ЍE�P�0 ����M�Q�@�@�ЋM����G��^�E�P�u ��_[��]Ë����  ��t5���V�u��@\�@,�Ѓ���u�M��r �M�V�q �E�   �u���u�M��^�  ���}���������E���t�����M�Q�@�@�С���M�Wj�h���@Q�@�ЍE�P��/ ����M�Q�@�@�Ѓ����u��Y| ���y WV����| �E�^P�/t ��_[��]�������U��SVW�}���u�' ���^����   �N0����   ���Q�@�@�Ѓ�����   �����  ����   ���S�@@�@,�Ћ�����؋Q��j h�  ���   �҅�tm�����j h�  �@�@0�ЋN0�-_ �N0j jjZjZ��_ �N0j j j �` Wh�  ���N ��t j ����G ��tj jh   �v0���` _^[]� �������U���u��j h&� �[� ]� �������U��V�u��j h�� �:� ����tj j h�� ��1 ����^]� ������������U���V���W��f/��E��E��$v�% ���# �]��E�������FW�f/��E��E��$v��$ ��# �]��E����F���FW�f/��E��E��$v�$ ��q# �]��E����F���FW�f/��E��E��$v�`$ ��9# �]��E����F^��]�����U���@SVW����$ �؅�t7���h-� S�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3����z ����M�Q�@�@�С���M�j j�h,��@Q�@�С���M�Q�@�@�ЋE��HK������  �$����������  j ���.h���s  ���k���g  ���6����[  �vP����  �L  j �vP�������;  ��������/  S�vP��誋���  �FH�E�jP���E��n��������o ��E��X���1�FH�E�jP���E��;��������o ��E��\���vP�N ���$�  �   ����s ���+�����P��s �NP�+�����P���  j�E���P����������o �vP��N ������$�^  �F�vP����������t6�
��$    �I ���j hȴ ���   �ϋ@���vP�����  ����u֋�� ����M�Q�@�@�С���M�j j�h8��@Q�@�С���M�Q�@�@�Ѓ���j ��q _^[��]� ��́ف��Z�����Z�Z�Z�+�;�n�݂��Z������U��W�}��t)VW��������tj j j���k�  W���#�  ����u�^_]� �������U��Q���SVW�@@�}j W�@8�M��Ѓ���3����V�R\��t'V�����  ����tjj j����  �M�W�����}F��c|�_^[��]� ����������U���   W���P ��  �GHW��oW(S�E��oG8��h���f(��\O0�\��,��,؉E���  �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3�V�wP���U���������OTj h[  �R���   �҉E���L  �O V�E�P�����E���h����Y����P�E��E��Y���E��^�  �U��u��_h��\M��@�\E��}��Y��Y��Y��u��M��Oxf/��E��Y�vf(��f(�f/�v�]���M��W`�Gpf/�vf(��f(�f/�v�U���E�f/�w(�f/�w(Ѓ}� �E��\e��\m�fn�����\�fn�����\��E�tO�X�f/��   �X�f/���   �E��X�f/���   �X�f/���   3�9Ej ��Pj��   �E��E��u��M��E��E��E��E��f/��E���   �X�f/�v{�E�f/�rp�X�f/�vf�E��XE��X}��E��u��M��}��E��E��E��f/��E�r&f/�v �E�f/�rf/�v3�9Ej ��Pj�jjj �����  �wP����  ���O �������^[_��]� ��������U��IW�}��t4���V���   �@X�Ћ���t3���;���P�L�  ����  ����u�^�} tj Wh�� �) ��_]� ���U����  ����u�M�@@�@,�ЋM���E�j �d� �8�  �P  ����M�Q�@�@�С���M�j j�hx��@Q�@�С���u���   �@8��H������  �$�Ԏj h��������D������M�Q�����Q�@�@�Ѝ�����  j hĻ�������������M�Q������Q�@�@�Ѝ������V  j h̻�M���������M�Q�M�Q�@�@�ЍM��*  j hػ��H����������M�Q��H���Q�@�@�Ѝ�H�����  j h��M��|������M�Q�M�Q�@�@�ЍM���  j h��������M������M�Q������Q�@�@�Ѝ������  j h ���h����������M�Q��h���Q�@�@�Ѝ�h����_  j h���h�����������M�Q��h���Q�@�@�Ѝ�h����*  j h���H����������M�Q��H���Q�@�@�Ѝ�H�����  j h��������y������M�Q������Q�@�@�Ѝ�������  j h,���(����D������M�Q��(���Q�@�@�Ѝ�(����  j h<���(����������M�Q��(���Q�@�@�Ѝ�(����V  j hD��M���������M�Q�M�Q�@�@�ЍM��*  j hP��������������M�Q������Q�@�@�Ѝ�������  j h\��M��|������M�Q�M�Q�@�@�ЍM���  j hh��M��P������M�Q�M�Q�@�@�ЍM��  j hx��M��$������M�Q�M�Q�@�@�ЍM��q  j h����x�����������M�Q��x���Q�@�@�Ѝ�x����<  j h����X�����������M�Q��X���Q�@�@�Ѝ�X����  j h����8����������M�Q��8���Q�@�@�Ѝ�8�����  j h��������V������M�Q�����Q�@�@�Ѝ�����  j h���������!������M�Q������Q�@�@�Ѝ������h  j h����������
������M�Q������Q�@�@�Ѝ������3  j h���������
������M�Q������Q�@�@�Ѝ�������   j h̼�������
������M�Q������Q�@�@�Ѝ�������   j hԼ��x����M
������M�Q��x���Q�@�@�Ѝ�x����   j h���X����
������M�Q��X���Q�@�@�Ѝ�X����bj h���8�����	������M�Q��8���Q�@�@�Ѝ�8����0j h��������	������M�Q�����Q�@�@�Ѝ�������Q�@�@�Ѓ�����M�Q�M�h<  �@�@8�С���M�Q�@�@�Ѓ��u�M��u�u�u��  ��]� �����$�P�������P������$�P�����݋	�>�s���݌�G�|�����J�������������������������U���X���SVW�@@�u�M��@,�Ћ]�����ˉ}�j �0� �8�  �z  ����u���   �@8�Ћ�������Q��j h�  ���   �ҋ�����E�P�I�I�ы��j j�h���A�M�Q�@�ЋM��E���VP�����������E�P�I�I�ы���A�M�QV�@�С���M؃��@�@<�Ћ��j�j��Q�M�QP�M؋BL�ЋM��E�WP�r���������E�P�I�I�ы���A�M�@Q�M�Q�С���M���@�@<�Ћ��j�j�V�Q�M�P�BL�С���M�Q�M�h<  �@�@8�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�ЍM���   j ��衆 �8�  �	  �����j h�  �@���   �Ћ�����u���   �I8�ы�����E�P�I�I�ы��j j�h���A�M�Q�@�ЋM��E��VP�G����M�P�E�PW�E�P�5���P�E�P������P�E�P����������Q�M�Ph<  �B8�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�ЍM���Q�@�@�С���M�Q�@�@�Ѓ��u�M��uS�u�
�  _^[��]� �U���   ����u�M�@@�@,�ЋM���E�j �D� �8�  ��  ����M�Q�@�@�С���M�j j�hx��@Q�@�С���u���   �@8�Ѓ����  �$���j hT���x����%������M�Q��x���Q�@�@�Ѝ�x����2  j hd��M���������M�Q�M�Q�@�@�ЍM��  j ht��M���������M�Q�M�Q�@�@�ЍM���   j h���M��������M�Q�M�Q�@�@�ЍM��   j h���M��o������M�Q�M�Q�@�@�ЍM��   j h���M��C������M�Q�M�Q�@�@�ЍM��Yj h���M��������M�Q�M�Q�@�@�ЍM��0j h����h�����������M�Q��h���Q�@�@�Ѝ�h������Q�@�@�Ѓ�����M�Q�M�h<  �@�@8�С���M�Q�@�@�Ѓ��u�M��u�u�u��  ��]� ْ�:�f���������������U���x����u�M��@@�@,�ЋM���E�j �ׂ �8�  ��  ����M�Q�@�@�С���M�j j�hx��@Q�@�С���u���   �@8�Ѓ����  �$���j h���M��������M�Q�M�Q�@�@�ЍM���   j h���M��������M�Q�M�Q�@�@�ЍM��   j h̻�M��c������M�Q�M�Q�@�@�ЍM��yj h���M��:������M�Q�M�Q�@�@�ЍM��Pj h���M��������M�Q�M�Q�@�@�ЍM��'j hĽ�M���������M�Q�M�Q�@�@�ЍM����Q�@�@�Ѓ�����M�Q�M�h<  �@�@8�С���M�Q�@�@�Ѓ��u�M��u�u�u��  ��]� F�r���Ǖ��U���H���V�u�M��@@�@,�ЋM���E�j �� �u�8�  �,  ����M�Q�@�@�С���M�j j�hx��@Q�@�С��V���   �@8�Ћ��P�E�P�I�A(�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M��<�@�@<�Ћ��j�j��Q�M�QP�M�BL�С���M�Q�@�M��@8h<  �С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ћu���u�M�V�u�u�)�  ^��]� ��U����V�uW���   ���FP�B<��3����_8�>���G@�   _^]� ������U���@���@�Mf/�VW��w���f/�v(�(��^F(f.���E���D�T  �}�E�P���N(��  �E���P��  �m�W��M��E��u�}f(��\]��f(��\U�f.��E��E��E�W��fE���D{	�^��]��E�f.ğ��D{	�^��U��Ef.ğ��DzW�fE��U��]���]��U��^��^��m��M��E��f.��E��E��E��E���Dzf.ğ��DzW�fE��U��]���Y��Y��\���\��ċ�f��0��  �F(�����$�G�  W���/,��_^��]� �������U��S�]V��9^P��   W�� �ȅ�t7���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ����3�S�N �^P�+���FP��t1jP���;���j j hɴ �= j �vPh�� �. ��_^[]� j j h�� � ��_^[]� ������������U���P���W�VW�����@�$�O ���   j	�С���O ��W��]��@�$j���   �С���O ��W��]؋@�$j���   �С���O j j�]�@���   ��j j���E��  W��E�    ���ύE�$V�E��� �D$�E��D$�E��D$�E�$P�l ����M�Q�@�@�С���M�j j�hx��@Q�@�Ѓ���rgdft{��tcpf��   ����M��E�YX�Q�@�E�@�С���M�j j�hг�@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�ЍM��u�E�M��Yh����Q�^��@�@�E�С���M�j j�h̳�@Q�@�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�ЍM���Q�@�@�Ѓ�����M��Ej0j �@j	j����@$�$Q�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@���E��,W�f.����D����@zQ�@�M�Q�С���M�j j�h|��@Q�@�С���M�Q�M�Q�@�@�С���M�Q�@�@�Ѓ� ��   �@<�M��Ѝp���~!���V�A�M�Q�@4�Ѓ�f��0uN��ߡ���M�VQ�@�@4�Ѓ�f��.uN����M��P�FPj �E�P�BP�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M�Q�@�@�Ѓ�����M��E�  �E    Q�@�@�С���M�Q�M�Q�@�@�С���MЃ��@�@<�Ћ��j�j��Q�M�QP�MЋBL��j j �EЋ�P�EP�n ����M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ�_^��]� ��U���TSVW���}�� �ȉM���t8���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E���E�    ������j j �@�@�Ћ؋�j�E��]�P������} �.  ���3�������   �@X�ЋЅ��  ���F���   �ʋ@(�ЋЅ�u����   ����M�Q�@�@�С���M�j j�hx��@Q�@�С���M��E�    �E�    Q���   �M�Q�@$�С���M����@Qj �ˋ��   �С���M�Q���   � �С���M�Q�@�@�С���M�Q�@�@�С���M�j j�h���@Q�@�С���MЃ��@Qh�� �ˋ@8�С���M�Q�@�@�Ѓ��Gj j
S�u�u�p计 �u���؉]��t����+ V��  ������  ����M�Q�@�@�С���M����@QS�M����   Q����Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M�Q�@�@�С��������P��'  j P���   �Ѓ} �Euj�E���P�Ӱ���o ��oE��M��E���� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ��M��T* �E�Phacpihbyek�1� ����M����@j haqpi���   �ЍM����z* ��u�M�V蜭���M�P�ci���E3�=�� uSSP�/ ���/  =�	 ��   �oE������u�� ���jj ���@��V�@�С���M�VQ�@�@�ЋM���h�� �  �؅���   ���S�@@�@,�ЋM��Q�ϵ ����������   ��j V���   �ҋ��Vh�  �A�ϋ@p�С��j S�@@�@8�Ѓ��ȋj �Rh�e�M��-�� t+��&t����Q�:h�� ���XV���؅�u:����hմ �hG  ���:V���؅�u����h�� �oE���� �:X���؋u����   ���~   ���j S�@@�@8�Ѓ����} t.���j �R\��tj�u��j �ߴ  ����PT��t=jS�u�.�E��cu"3������V�P\��uF��c|��j�u��V�jSP��藴  �M�j �Q �M��� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�С���M�Q�@�@�ЋE��_^[��]� _^��[��]� ��������������U���@VW�M���  ���M��u��' ��u�M������' ��_^��]� ���Sh-� V�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��E����3ۉ]��K��u3��������   �@X�Ћ�����M�Q�@�@�С���M�j j�h���@Q�@�С���M���@Qh�� �M��@8�С���M�Q�@�@�С���M�Q�@�@�С���M�j j�hx��@Q�@�С���M��E�    �E�    Q���   �M�Q�@$�С���M�� �@Qj �M����   �С���M�Q���   � �С���M�Q�@�@�Ѓ����  ��� �d$ ���9�  ������E�P�I�I�ы����j �x����DIj�P�E�P�A�Ѓ������  ������E�P�I�I�ы���A�M�QV�@�С���M���@�@<�Ћ��j�j��Q�M�QP�M�BL�С���M��P�E�P������P�B8�С���M�Q�@�@�С���M�Q�@�@�С�����@WS�@p�M��Ћ���  ��C��������]��u�E��M�j j
Q�u�@�u�p�� ������~R���� u�M����[�M��)% ��_^��]� ����M�j V�P��'  P�Bl�Ћ���jV������M�V����[�M���$ ��_^��]� �������������U���E�3� �E� �E�"� �E� ]����������V���vP�N ����j ���)M ^� �����U�������E�� �$�$��]��3���������������U���0VW��M�hTCAb��# �M���# ���M ���Phdiem�Q�M�B4�С���M�j havem�@�@4�ЍE��E�    P�vX���E�    hsuom�N ����M�j hxvpi�@���   �ЉE��MС��j hyvpi�@���   �ЉE��΍E�P�E�P��T ����M�j haqpi�@���   �Ћ����j havpi�Q�MЋ��   �҅���   ����M�j hrdem�@�@4�ЍE��P�qL fnM���fnE���P�ǋ΃���P���W�����vX���f���H7��j ���K j �� ���FX    ��j ��L �dfnM���fnE���P�ǋ΃���P���W�����vX���f���*4��j ���1K ����M�jhrdem�@�@4�ЍE��P�K �M��g" �M��_" _^��]� ������������� ��������VW���7� �ȅ�t5���h-� Q�@L���   �ЋЃ���t���j R�A@�@8�Ѓ��3��wP��萸������t1j ��豩  ��t���V�  �؋��@P�	�  �wP����  ����u�j ���PJ _^��������������U��W�u���O�# �u�O�# �   _]� ����������U���HS�]���E�VW��u膤���؅�u3��  脷���u�E��( ��������  ���S����@V�@�С���MVQ�@�@�Ћu��E؃���P�  ����ЋA�MQR�@�С���M�Q�@�@�Ѓ��E��P�1�  S���	�  ���W��Mj hM  �@fE؋��   �Ѓ� ��   Ht����   E(E��   �Eȋ�P���  ����Y���M��H�E��Y��P�M���  �E��X �E��@�XE��E��E��E��E��E��E��E��E��E��%W�(��M���U�E�(�����E��M��oE؃��ϋ�� 諭  �}  tjj j���8�  ����NW���   �@h�ЋM$��tGWj,�� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ѓ�����EP�I�I�у���_^[��]�0 ������U����} SVW��t5�K��t.������   �@X�Ћ���t��j ���7�  ����  ����u�h*� �`& ��������   �������IV�I�ѡ���MVQ�@�@�Ѓ��E���P��  ����ЋA�MQR�@�С���M�Q�@�@�Ѓ��E��P��  �} t	j����  ����KW���   �@h��j Wh�� � ����MQ�@�@�Ѓ���_^[��]� ������������U��E��x;A,}�E��x;A0}	�   ]� 3�]� ������U��V�u���r�  �N<��t�x �F<    ^]� ����������U��]�G�  �������U��V�u���2�  �N4��t����@ �@T���F4    ^]� ��U���SV��N��t:������   �@X�Ћ؉]���t!��    �����  ��u#����  �؉E���u�E^[� ����3���]� ��t�WS��3��#����؅�tU���j S�A@�@8�Ѓ��E�3��d$ ���V�R\��tV���,�  ;Eu;}t.G�E�F��c|��u����~�  �؅�u��E_^[� ����3���]� �E_�0��^[��]� ����U�����W��Mf(��\}L���   f(�f(ύI �t�Y���t
f(��Y���f(ϸ   f(�t�Y���t
f(��Y����ML�   f(�t�Y���t
f(��Y����ML�   f(���I �t�Y���t
f(��Y����ML�   �Y ��Ym�YU<�M�f(��Y ��M��M��E��Y��Y��YM�YE,�X�f(��X��X��	f(ύd$ �t�Y���t
f(��Y���   f(㐨t�Y���t
f(��Y����uL�   f(�f(Өt�Y���t
f(��Y���   �t�Y���t
f(��Y����E����M��Ym�Y]D�Y��Y��YE$�YM4�X��X��X��A��]�L �������̋IV3���t"������   �@X�Ѕ�t����F��  ��u��^�U���`SVW�u���������������W�@�@�С���MWQ�@�@�Ѓ��E���P�؜  ����ЋA�MQR�@�С���M�Q�@�@�С���]S�@�@�С���MSQ�@�@�Ѓ��E   ��I ��tj���u�  ������E�P�I�I�ы���A�M�QW�@�С���MЃ��@S�@x�Ѕ�tD�u��輟  ���MС��Q�@�@�Ѓ���u�����EP�I�I�у���_^[��]� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M��uQ�@�@(�Ћ�����E�P�I�I�ы���A�M�QW�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�MQ�@�@�С���M���8�@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�С���M��@�@Q�M�Q�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�SQ�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M��EQ�@�@�Ѓ���������U���`S��VW�K��u3��������   �@X�Ћ��������@W�@�С���MWQ�@�@�Ѓ��E���P��  ����ЋA�MQR�@�С���M�Q�@�@�С���]S�@�@�С���MSQ�@�@�Ѓ��E   ����tg����  ������E�P�I�I�ы���A�M�QW�@�С���MЃ��@S�@x�Ѕ�tA���?�  ���MС��Q�@�@�Ѓ���u�����EP�I�I�у���_^[��]� ����M�Q�@�@�С���M�j j�h���@Q�@�С���M��uQ�@�@(�Ћ�����E�P�I�I�ы���A�M�QW�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�MQ�@�@�С���M���8�@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�Q�@�@�С���M��@�@Q�M�Q�С���M����@�@<�Ћ��j�j��Q�M�QP�M��BL�С���M�SQ�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���M��EQ�@�@�Ѓ������������U��V�uW�u���uV��  ���V�@@�@,�Ћ�������Q��jh�  ���   ��������G4����$h�  �A�΋��   ���_8_3�^]� �������U��V�uW�u���uV蚯  ���V�@@�@,�Ћ�������Q�$�A��h�  ���   ��������_8������$h�  �@���   ���_@�����jh�  �@���   �ЉGH�Ρ��j h�  �@���   ��������GL�Ρ���$h�  �@���   ���_P�����jh�  �@���   �ЉGX�Ρ��jh�  �@���   �ЉG\3�9GHt
�G8�G@_^]� ������U���0V�uW�u���uV�g�  ���V�@@�@,�Ћ�������Q��jh�  ���   �҉Gh�M���W�QfE�M��E��@h�  Q�΋��   ��jh�  ���o �G8�~@f�GH����@���   ��(��M�Gl���fE�Q����M��E��@h�  Q�΋��   �Ѓ����o �GP�~@f�G`�������$h�  �@���   ���_p_3�^��]� �������������U���0W�u���u�u�9�  ����u�@@�@,�Ћ����W���fE��E��A�M�Qh�  �MЋ��   Q�����o �G8�~@3�f�GH_��]� �����������U��V�uW�u���uV躬  ���V�@@�@,�Ћ�������Q��jh�  ���   �҉G4���j h�  �A�΋��   ��h!D h�  �ΉG8�� �G<_^��t�u���k ��t3�]� �����]� ������U��V�uW�u���uV��  ���V�@@�@,�Ћ�������Q��j h�  ���   �҉G4���j h�  �A�΋��   �ЉG83�_^]� �����U��S�]VW�u���uS詫  ���S�@@�@,�Ѓ��E�G4    �   V��著  ��t�w4F��
~����]��jh�  �@���   �ЉG8�����W����$�@h�  ���   ���_@�����jh�  �@���   ��h�e h�  �ˉGH� �GL3�_^[]� �������U��V�uW�u���uV�ڪ  ���V�@@�@,�Ћ�������Q��jh�  ���   �҉G4���jh�  �A�΋��   �ЉG8�Ρ��jh�  �@���   �ЉG<�Ρ��j h�  �@���   �ЉG@�Ρ��jh�  �@���   �ЉGD�Ρ��jh�  �@���   �ЉGH3�_^]� �����U��V�uW�u���uV���  ���V�@@�@,�Ѓ�����h�e h�  �f ������G4����$h�  �A�΋��   ���_8_3�^]� U��V�uW�u���uV芩  ���V�@@�@,�Ћ�����0�Q�$�Q��h�  ���   ��������_8������$h�  �@���   ���_@�����jh�  �@���   �ЉGP�Ρ��jh�  �@���   �ЉGT�Ρ��jh�  �@���   ��h�f h�  �ΉGX�R �G\��tk��蔈 ��~`�O\3�膈 ��~R������ϋ��   �@T�ЋO\VP脇 ��u#�O\V�� ��t#���jW�@H���   �Ѓ��O\F�4� ;�|�_3�^]� ��������U��V�uW�u���uV�*�  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ���_8�����W��΋@�$h�  ���   ���_@�����j h�  �@���   ��������GH�Ρ���$h�  �@���   ���_P�����jh�  �@���   �ЉGX3�_^]� ��U��S�]VW�u���uS�I�  ���S�@@�@,�Ћ�����x�Q�$�Q��h�  ���   ���_8�����jh�  �@���   ��h�f h�  �ΉG@�s �GD��tl��赆 ��~a�OD3�视 ��~S�I ����ˋ��   �@T�ЋODVP褅 ��u#�ODV�7� ��t#���jW�@H���   �Ѓ��ODF�T� ;�|�_^3�[]� �������U��V�uW�u���uV�J�  ���V�@@�@,�Ћ��W�Q���$h�  �Q�΋��   ���_8�����W��΋@�$h�  ���   ��������_@������$h�  �@���   ��������_H������$h�  �@���   ��������_P������$h�  �@���   ��������_X������$h�  �@���   ���_`_3�^]� �U��V�uW�u���uV�*�  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ���_8�����j h�  �@���   �ЉG@3�_^]� �������������U��V�uW�u���uV誤  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ��������_8������$h�  �@���   ���_@�����W��΋@�$h�  ���   ���_H�����jh�  �@���   �ЉGP3�_^]� ��������������U��V�uW�u���uV�ڣ  ���V�@@�@,�Ћ��W�Q���$h�  �Q�΋��   ���_8�����W��΋@�$h�  ���   ���_@�����W��΋@�$h�  ���   ���_H�����j h�  �@���   �ЉGP�����W����$�@h�  ���   ���_X�����W��΋@�$h�  ���   ���_`�����W��΋@�$h�  ���   ��������_h������$h�  �@���   ���_p�����j h�  �@���   ��������Gx�Ρ���$h�  �@���   ��ݟ�   _3�^]� ������U��V�uW�u���uV�:�  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ���_8�����jh�  �@���   �ЉG@3�_^]� �������������U��V�uW�u���uV躡  ���V�@@�@,�Ћ�������Q��j h�  ���   �҉G4���jh�  �A�΋��   �ЉG8�Ρ��j h�  �@���   �ЉG<�����W����$�@h�  ���   ��������_@������$h�  �@���   ���_H�����W��΋@�$h�  ���   ��������_P������$h�  �@���   ���_X����@��������   ���$h�  ���_`�����W��΋@�$h�  ���   ��������_h������$h�  �@���   ��������_p������$h�  �@���   ��������_x������$h�  �@���   �������ݟ�   ������$h�  �@���   ��ݟ�   _3�^]� ��������������U��V�uW�u���uV芟  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ���_8�����W��΋@�$h�  ���   ���Z� �G@�Ρ��jh�  �@���   �ЉGD3�_^]� ���U��V�uW�u���uV��  ���V�@@�@,�Ћ�������Q��j h�  ���   �҉G4���j h�  �A�΋��   �ЉG8�����W����$�@h�  ���   ��������_@������$h�  �@���   ���_H�����jh�  �@���   �ЉGP3�_^]� ����������U��]��  �������U��V�uW�u���uV���  ���V�@@�@,�Ћ�������Q��j h�  ���   ��������G4����$h�  �A�΋��   ���_8_3�^]� �������U��SV�uW�u���uV�y�  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ���_8�����W��ˋ@�$h�  ���   ���_@�����jh�  �@���   �ЉGH3���L�����j �P��M  P���   ��F����|�_^3�[]� �����������U��V�uW�u���uV誜  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ��������_8������$h�  �@���   ���_@�����j h�  �@���   �ЉGH3�_^]� ���U���u�u�u��  3�]� ���������U���0V�uW�u���uV��  ���V�@@�@,�Ћ�������Q��j h�  ���   �҉G4���jh�  �A�΋��   �ЉG8�Ρ��j h�  �@���   �ЉG<�����W����$�@h�  ���   ���_@�����W��΋@�$h�  ���   ��������_H������$h�  �@���   ��������_P������$h�  �@���   ��W��_XfE����M�Q�E��M�h�  �@Q�΋��   �ЍM�Qh�  �o �M�Q�G`���~@f�Gp( ����fE��X��E��@���   �ЍM�Qh�  �o �M�Q�Gx���~@fև�   W����fE��E��@���   ��jh�  ���o ���   �~@fև�   ����@���   �Љ��   3�_^��]� �����U��V�uW�u���uV�ʙ  ���V�@@�@,�Ћ�������Q��j h�  ���   �҉G4�����W��$�A��h�  ���   ��������_8������$h�  �@���   ���_@�����jh�  �@���   �ЉGH�Ρ��jh�  �@���   ��h�e h�  �ΉGL��  �GP3�_^]� ������U��V�uW�u���uV�ژ  ���V�@@�@,�Ћ�������Q�$�Q��h�  ���   ���_8�����jh�  �@���   �ЉG@�Ρ��jh�  �@���   �ЉGD�Ρ��jh�  �@���   ��h�f h�  �ΉGH���  �GL��tu���x ��~j�OL3�� x ��~\�
��$    �I ����ϋ��   �@T�ЋOLVP��v ��u#�OLV�w ��t#���jW�@H���   �Ѓ��OLF�w ;�|�_3�^]� ��������U��V�uW�u���uV蚗  ���V�@@�@,�Ћ�������Q��j h�  ���   �҉G4���jh�  �A�΋��   �ЉG8�Ρ��jh�  �@���   �ЉG<3�_^]� ���������U��V�uW�u���uV�
�  ���V�@@�@,�Ћ�����0�Q�$�Q��h�  ���   ��������_8������$h�  �@���   ���_@�����W��΋@�$h�  ���   ���_H�����jh�  �@���   �ЉGP�Ρ��jh�  �@���   �ЉGT�Ρ��jh�  �@���   ��h�f h�  �ΉGX��  �G\��ti����u ��~^�O\3���u ��~P����ϋ��   �@T�ЋO\VP��t ��u#�O\V�tu ��t#���jW�@H���   �Ѓ��O\F�u ;�|�_3�^]� �����U��W�u���u�u茕  ����u�@@�@,�Ћ�����ЋA��j h�  ���   �ЉG43�_]� ���U��SVW�u�}���uW�9�  ���W�@@�@,�Ћ�����ϋ����   �RT�ҋ��hK  Ph�  �Q�΋Bl��h.� P�C4�zp������t_^�����[]� �K4��t����u�@ �@P��_^[]� _^3�[]� U��V�uW�u���uV蚔  ���V�@@�@,�Ћ�������Q��j h�  ���   ��j h�  ��fn�����G8����@���   �Ѓ���fn�����G@W�����$h�  �@���   ���_H�����W��΋@�$h�  ���   ���_P�����W��΋@�$h�  ���   ��������_X������$h�  �@���   ��������_`����$h�  �@���   ����������_h������$h�  �@���   ��������_p������$h�  �@���   ���_x_3�^]� �����������U��} SW�}��tM�K��t6���V���   �@X�Ћ���t��3���;���P���  ���
�  ����u�^j Wh�� �6� ������KW���   �@h��_[]� ��������̋A�������������U����}u{V�u��    tm�E��E�  P�E��E�    P�E��P�E�P�E�P��W ��u�����ȉE��M��M��E��M��P�E�P�J �M�E�j j�j QP���   �����^��]������U��}uj h�� �� ��]�������U����}u|V�u�E�P�E��E�  P�E�E�    P�E���P�E�P�'W ��u�����ȉE�Q�M���   P����^��]ËM��E��M��P�E�P��I �M�E�QP���   �����^��]�����U���   VW��� t�u�u�u�uV軒  ��_^��]� �u��j �}  j�ΉE�	}  j�Ή�t�����|  �MW��E�W�f(������x������E�fM�fM�fM�fM���tL���j Q�@@�@8�Ѓ��M���u�u�uQ�ȋBH����x���W��o fE�fE��~@�E���t�����tG���j Q�@@�@8�Ѓ��M���u�u��t���Q�ȋBH���o�~hfM�fM���x���� ��   ����   ���j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$�,��M��%�M���M���M��XM��XM��Yh�W��M�f/�v
(��M�����f/�v(��M���M����� ��x���t�\�(��M�fMЋG4W�HfEȃ��i  �$�<�fE��]��E�f��M  �E�f/�vf(��f(��M��u�f/�w(��E��}�f/�w(�f��E��  �}�f(��u�f(��YM�(��YE��Ye�f��M���  fE����]��ă��f�h��� f�X�E�P�P���o ��4�~`�E��  fE����]��ă��f�h��� f�X�E�P�JQ���fE����]��ă��f�h��� f�X�E�P�Q����E�f/�vf(��f(��U��M�f/�w(��E��}�f/�w(�f��E���  fE����]��ă��f�h��� f�X�E�P�/R������fE����]��ă��f�h��� f�X�E�P�R��������}�f(��u�f(��XM��Xe�(��XE�f��M��R  fE����]��ă��f�h��� f�X�E�P�5S���q���fE����]��ă��f�h��� f�X�E�P��S���=���fE����]��ă��f�h��� f�X�E�P�=U���	���fE����]��ă�� f�X���f�h�E�P�iS�������fE����]��ă��f�h��� f�X�E�P�EW������fE����]��ă��f�h��� f�X�E�P��X���m���fE����]��ă��f�h��� f�X�E�P��Y���9���fE����]��ă��f�h��� f�X�E�P��Z�������U��}��M��\��u��@��\��e��\�fT�fT�f�fT��U��k  �E�f(��]�����X��u��Y�(��}��YE��\��E��X��Y��Y��\��E��X��Y�f��Y��]��\���  �}�f(��u�f(��\M��\e�(��\E�f��M���  fE����]��ă��f�h��� f�X�E�P��\�������fE����]��ă��f�h��� f�X�E�P�<]������fE����]��ă��f�h��� f�X�E�P�]������fE����]��ă��f�h��� f�X�E�P�T^���P���fE����]��ă��f�h��� f�X�E�P�]������fE����]��ă��f�h��� f�X�E�P�l^��������}�f(��u�f(��\U����f(��\M��\e��X��X��X�f��U��Q�}�f(��u�f(��XU����f(��XM��Xe��\��\��\�f��U��W��}��u��U��M��\���x����\��E��\�E�Y��Y��Y��G8�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� ����������?�W������H�y�����*�\�������,�`�������C������I�}������]�U������$  SVW��� t�u�u�u�uV�'�  ��_^[��]� �Mj �s  �M��j�\$�rs  ������L$��u�EW� �@_^[��]� � �]��   ����   ���j V�@@�@8�Ѓ��L$x��uSVQ���RH�GH��wx�$�P��T$x�6��$�   �+��$�   � ��$�   �XT$x�X�$�   �Yh����W�f/��T$v(��T$�"f/�v(��T$��T$W����� tf(��\�f(��T$�WۋGL�   �\$0W��\$8�щL$�T$f�$�   ;�wU�$�`��L$�T$�D�   �щL$�T$�3�   �щL$�T$�"�OX���L$%  �yH���@uA�L$�щL$�O8fn��������t$j V�@@�^ȋ@8fn�����L$x�O@�^��L$h�Ѓ��L$H��uSVQ���RH�O8W�f.��o �~X��\$h�d$x��$  ��Dz*�\ �   �t$�T$pt�E� f�X_^[��]� �t$�G@f.��Dz�D$   �T$`f.ʟ��Dz
f.��D{���$�   W�f�$�   f�$�   f�$�   f�$�   ��tjh��$�   SP��� ���L$����  ��$�   �A���$�   ��$�   ��$�   �\$`�+��d$ �����l$(�D$@fn�����Y��X���$�   ���  �L$�F��+L$D�������	��$    ����$�   �\Cfn�����Y��YT$p�X���$�   �\K��$�   �\�Y��Y��X��X�蜾 �G\f(ȃ� ��   H��   H�Q  �G8f/��B  �^ȡ��j �@@�@8����t$�\���$�   �Ѓ���$�   ��uQ�t$�L$TQ���RH��$�   �D$H�L$P�T$X�Y��Y��Y��XD$(�XL$ �X\$8�XT$0f(�f(��l$(�d$ �T$0�\$8�   �G8f/���   ���j �t$�@@�@8�Ѓ���$�   ��uQ�t$�L$TQ���RH�D$H�XD$(f(��D$P�XD$ �l$(f(��D$X�XD$0�d$ �D$0�D$8�X���D$8��d$ �l$(�F�L$D�"����\$`�t$�L$�D$@�S@I�D$@�L$������D$8W�f/�v(����^��t$h(�(��YL$0�Y��Y��+�oD$x�t$h��$�   ��$�   f���$�   �  ��$  u(Ճ$ ��$   u(܃( u(��D$�\��\܋E�\��Y��Y��Y��GP�X��X�_�X�^�\��\�[�\��Y��Y��Y��X��X��X�f��f�H��]� r�z�����F�P�a�r�U���PVW��� t�u�u�u�uV�n�  _��^��]� �MSj ��l  �M��j�l  W�W��E�������E�fM�fM���t=���j S�@@�@8�Ѓ��Mȋ�u�uSQ���RH�o fE�fE��~@�E�� [��   ����   ���j V�@@�@8�Ѓ��Mȋ�u�uVQ���RH�GH��wc�$����E��%�E���E���E��XE��XE��Yh�W��E�f/�v
(��E�����f/�v(��E���E����� t�\�(��E��h fE��m��u�f��E�tE�  t�_8f/�w�]ȃ$ �U�t�G@f/�v(Ѓ( t�GHf/�v(��
�U��]ȃl t<�  t�GPf/�v(؃$ t�GXf/�v(Ѓ( t�G`f/�v(��M��\��E��\��\�E�Y��Y��Y��Gp�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� �I `�g�n�u�����U��y t�u�u�u�u��  �E]� �oA8�E� �~AHf�@]� �����U���8VW��� t�u�u�u�uV�  ��_^��]� �Mj ��i  ��W�WɅ��_  ���j V�A@�@8�Ѓ��Mȋ�u�uVQ�ȋBH�ЋO4�Ѓ���~J�o�E�����   �$���o����� �~Bf�@�E�P�L5������{�o����� �~Bf�@�E�P�#5�����H�Q�o����� �~Bf�@�E�P��4�����H�'�M�� �M���E��XE��X��Yh�(ȋG8�M�Ht3HuB�E�����Ɯ ����]��E��\�fT@��\���E���蚜 �]��M��O<�Eȃ��$P�4< �o �~H�E_^� f�H��]� �I ���7�a�h���������������U���`VW��� t�u�u�u�uV�}  ��_^��]� �Mj �
h  ��W��E�W�fE���2  ���j V�@@�@8�Ѓ��MЋ�u�uVQ���RH�O4���ofE��~J�M�;O8��   ItPIt(Ium�o����� �~Bf�@�E�P�qS�����5�o����� �~Bf�@�E�P��4������E�P�E�P��� ���o fE��~H�M��G8Ht>HtHuV����� f�H�E�P�T�����,����� f�H�E�P��2������E�P�E�P胒 ���o fE��~H�E� f�H_^��]� �E_^�f�@��]� ����������U���xSVW��� t�u�u�u�uV�|  ��_^[��]� �4 W�W�u�E�f�@_^[��]� �]��j �Ef  ����u�EW�� f�@_^[��]� ���j V�@@�@8�Ѓ��MЋ�u�uVQ���RH�G8�������   �$����oEЃ���� �~E�f�@�E�P�1����� �   �oEЃ���� �~E�f�@�E�P�~1�����@�W�oEЃ���� �~E�f�@�E�P�S1�����@�,�E��%�E���E���E��XE��XE��Yh��OL�E����$P��@ ���W��Hf/�v(��	f/�v(ʋw4f(�f.�fn������^���Dz����   �E��   f.ʟ��Dz(��   3���~6���$    fnЍH���fn�����Y��Y�f/�rf/�w��;�|�W�E_^[� f�X��]� ���p�L$�D$�$�_.�������%���]��E��E���~��G@��f.�V���Dz:�d  ���������V�|���M���Q�MQV�M�Q���RH�o �~X�g���W��]�fE�f(��E�W�fE���c  �E��t4P�W|���M���Q�MQ�u�M�Q���RH�o �~Xfe��]���]�W��M�W�f/���   �o@�\�f.���D{�X���\��^�(����$��)�����]���u�H t�w4��e�f�]��AN��~<V���c  ����t.V�{�����M���u�uVQ���RH�o �E��~@�E��U��Y���M��\M��]��X���\]��Y��Y��XM��X]�f(��M��\M��Y��XM�f���������f(��\o@�\�f.П��Dz(���\��^ʃ��$��(���G4���]�;�u�H tj��e�f�]��AF;�<V���b  ����t.V�z�����M���u�uVQ���RH�o �E��~@�E��U�W��Y���M��\M��]��\]��X��Y��Y��XM��X]�f(��M��\M��Y��XM�f������I ���������������������U���0VW��� t�u�u�u�uV��v  _��^��]� �Mj�*a  ����u�EW�_^ �@��]� ���j V�@@�@8�Ѓ��M��u�uVQ���RH�Mj ��`  ����u�E�oE�_^� �~E�f�@��]� ���j V�@@�@8�Ѓ��MЋ�u�uVQ���RH�4 �M��U��E�t!�G@�� tHt
Hu�M���U���E�8 t!�GD�� tHt
Hu�M���U���E��< t�GH�� t)Ht!Ht�M��E�oE�_^� f�H��]� (���(����������������U���pVW��� t�u�u�u�uV�^u  _��^��]� �MSj �_  �M��j�_  ���W��M����E�fM�fM���t=���j S�@@�@8�Ѓ��M���u�uSQ���RH�o fE�fE��~@�E�� [��   ����   ���j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$� ��E��%�E���E���E��XE��XE��Yh�W��E�f/�v
(��E�����f/�v(��E���E����� t�\�(��E��  fE��E�t �E��E��O4���$P�: �@��E؃$ �E�t �E��E؋O4���$P��9 �@��E��( �E�t �E��E��O4���$P�9 �`��~e��oUȋE�u��m��\��]��M��\��E��\��Y��Y��Y��G8�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� m�t�{���U���(  VW���}�� t�u�u�u�uV��r  ��_^��]� �uW�W��~T ��  �Mj �]  (�������U��M�f�8�����tA���j R�A@�@8�Ѓ���������uV�u�Q�ȋBH���o ��8����~@�E��P W��NTfE��E��o��   �E��~��   f�E��o��   �������~��   fօ ����o��   ��P����~��   fօ`���u�o��   �E��~��   f�E�3�9��  Q��3�9WTD�3��E����}��@�@X���Mȃ��E����J  �M��E���W�vT�@�@T�Ћ����E��x\ t>������   �M�RT���wP�E��H\�wM �M�3�9QX��3Ƀ����;���  �vTW�j ���j�o��   ��@  ������~��   fօ���W�f�p����M�fE��M���(  ���   Q�u��@��P�����RQ��d  ������Q�M�Q�����Q�M�Q��p���QWV�Ћu��8���  ���  �E    �E�    �9 t$�E�P�EP�FT��0  Q�ڋ ���} ��  ���   W�W�f(�u}���W��VTfE��M�f� �����0����H�� ���P�E�P��(  ��P���P�E�P�����P���   ��P��`  ���$jj WR���oe���4�~]��   �E��YE��FT�U��YU��X��E��YE��X���  �Y�f/�rZ��8  f.����D{4fT@�fWP���h����c� f(���h����"� f(��f(�fT@�f(�f�}��� ���G@�D$� f�X�� ���P��*���G8��$�o�~X�Y]�f������������Y�p����Y�x����Y��Y��Y�W�f/�v(�f/�v(�f/�vf(��E��X��E��E��X��E��E��X��Eء���}��vTG�@�}��@X�Ѓ�;�������E��M��Y�8����Y�@���f(��E��YE�fыE_^�f�@��]� ���U����   VW��� t�u�u�u�uV��m  _��^��]� �u��j �%X  j�ΉE�X  ������M�E���u�EW�_^ �@��]� � ��   ����   ���j V�@@�@8�Ѓ��M܋�u�uVQ���RH�GH��wd�$�  �M��%�M���M���M��XM��XM��Yh�W��M�f/�v
(��M��f/��v����M���M�� �Mt����\�(��M��GH�   W�W��U�fE�;�w)�$�0 �   ��   ��wX��%  �yH���@uF�O8fn�f(����f.��^؟�]���Dz
�   �U����j Q�@@�@8�Ѓ��M���u�u�uQ�ȋBH���o ��|����~@�E�E�W���T���f����f�$���f�4���f�D�����tjhP�����P�T� ��3��E���)  �E��E��E��E��G@fWP�fn�����E��YM��M��� �YEċE�X ������E��ɒ �YEċEj �u�X@���������@@�@8�Ѓ��������uQ�u�M�Q���RH�E��XE�E�@�E�f(��E��XE��U�f(��E��]��XE�f(��e�;��/�����~Ofn�W����f.���D{����^�(��Y��Y��Y��f(�f(�f(���]��U��eԃ  ��|���uf(Ճ$ �M�uf(ك( �u�uf(��E��\��\ًE�\��Y��Y��Y��GP�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� ������������l�s�z�U������  ��3ĉ�$�  �ES�]V�uW���D$D� t�uSPV�i  �p  �CTW�WɅ��V  fD$x�D$p    f�$�   �D$l    f�$�   Ǆ$�       �$�   f�$  f�$   f�$0  f�$@  f�$P  f�$`  f�$p  f�$�  f�$�  f�$�  ��$�  ���   �T$0���   ���   (��Y��L$H(��Y��\$8�X�(��Y��X��á f(�W�f.џ��DzW��L$`fD$P�<����^��L$0�T$8�\$H�Y��Y��Y��L$X�T$`�\$P�D$PP�CT���   ��P��$�   P�Fz �KT�T$t����������$  �o��   R�T$4��$�   R�~��   ��$�   ��$H  ���D$D    ��$8  �D$@    ��$   �o�$�   fք$�   fք$`  fք$H  fք$0  �~�$�   fք$  fք$�  fք$�  fք$x  �G8��$   ��$�  ��$�  ��$h  �@�$RQ��$  �Ѓ���uW��f�F��   �|$4�t�D tP�D$h�D$8��tD���    t;����L$D���   �@T�ЋL$8���   �ODP��B 3�9W@��3Ƀ����;�t��CT���   ���   �\�$�   �\T$x���   �\�$�   �Y��Y��Y��X��X��|� �^G8���W��\�f/�w(�f(�f��f�N��$�  ��_^[3��F� ��]� �����U����   VW��� t�u�u�u�uV��e  _��^��]� �u��Sj �$P  j�΋��P  j�ΉE�P  ����E��E����  ���j S�A@�@8�Ћu�M�����uVSQ���RH�M�~H�M��o �E�����  ���j Q�@@�@8�Ѓ��MЋ�uV�uQ���RH� �o �E��~@f�E���   �E����   P��g���M����uVQ�M�Q���RH�GH��wc�$���E��%�E���E���E��XE��XE��Yh�W��E�f/�v
(��E�����f/�v(��E���E����� t�\�(��E��WHW��_PW���X����^��^��U��]�f����f�(���f�8���f�H�����tjh�����VP�w� �U����]�W��%��f.џ��Dz
������'�E��\��^��YGX�X�����\G8�����f.ٟ��Dz
�� ����'�E��\��^��YGX�X� ����XG@�� ������j S�@@�@8�Ѓ��������uQS�M�Q���RH�  �u�uf(���M��$ �e�uf(���]��( �m�uf(���U��E��\��\܋E�\�[�Y��Y��Y��G`�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�P��]� �E[_^� f�H��]� �EW�[_^ �@��]� �I 9@GN����U������L  �y SVW�L$@t�u�u�u�uV�b  ��_^[��]� �Mj �pL  W�Wɋ��L$ �L$p�L$0fD$`fD$HfD$`��u�E�H_^[��]� �M��$�   f�$�   f�$�   f�$�   ��tjhQ��$�   P�� �M���D$P����\$`�D$(�D$H�D$H�D$h�T$D�D$8�\$�d$ �D$@�4�    fn������Y@8�XA��$�   ��$    fn�����Y@8�@@�X�D$x�� ��  H�  H�  9����   ���j S�@@�@8��fn����$�   �������u�D$QS�L$lQ���RH�\$�H�P� �Y��Y��Y��XL$(�XT$ �\$�XD$H�L$((��L$ �D$H��0� �p  ���j S�@@�@8��fn�0���$�   �������u�D$QS��$4  Q���RH�\$f(��Y �H�P�Y��XD$�Y�f(���  ��ı ��   ���j S�@@�@8��fn�ı��$�   �������u�D$QS��$L  Q���RH�\$� �H�P�Y��Y��Y��XD$H�XL$(�\$�XT$ �D$H�L$(�T$ ��� �]  ���j S�@@�@8��fn����$�   ���uQ��$�   ��   ��|� ��   ���j S�@@�@8��fn�|���$�   �������u�D$QS��$  Q���RH�\$f(��H�P�Y �Y��Y��XD$H�XL$(�\$�XT$ �D$H�L$(�T$ ���� ��   ���j S�@@�@8��fn�����$�   ���uQ��$  ����SQ���D$ �RH�\$� �H�P�Y��Y��Y��XD$(��XL$8�XT$0�\$�L$8�T$0�D$@G�M����������T$DB�T$D���f����D$H�Y��Y��X��ϖ �L$(�D$H�D$8�Y��Y��X�謖 �L$0�D$�D$ �Y��Y��X�(�膖 fT$H�E�L$_f�^�[f�@��]� �U����   VW��� t�u�u�u�uV��\  _��^��]� �MSj �VG  �M��j�JG  ������E�����  ���j S�A@�@8�Ѓ��M���u�uSQ���RH�o �E��E��~@�E�E�W���h���f�(���f�8���f�H���f�X�����tjhP��(���P�Ԙ ���GH觓 �YG@�X�(�����(����GH舃 �YG@���j S�X�0�����0����@@�@8�Ѓ���(�����uQS�M�Q���RH� �o �E��~@�E���   ����   ���j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$���E��%�E���E���E��XE��XE��Yh����W�f/��E�v
(��E�� f/�v(��E�����W��E�� t�\�(��E��W�  �oE��}��u�f��E�t$�P tf(��f(��M��\��YO8�X���M��$ �m�t$�P tf(��f(��U��\��YW8�X���U�( t�P t(��]��\��Y_8�X��E��\΋E�\��\�[_�Y�^�Y��Y��X��X��X�f��f�X��]� �EW�[_^ �@��]� ������������U���   VW��� t�u�u�u�uV��Y  ��_^��]� �u��j �%D  j�ΉE�D  ������M�E�W����  ���j Q�@@�@8�Ѓ��M���u�u�uQ�ȋBH�Ѓ �o �~H�E��E��M���   ����   ���j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$��M��%�M���M���M��XM��XM��Yh�W��M�f/�v
(��M�����f/�v(��M���M����� t�\�(��M��oE��E�P�EȍE��E�Pf�E��xn �G8���P �^(�t�E��G@�E��M�XE��E��E����v �E�W��O@�Y���Y���]��X���\��Y��X��M��E�P�E�P�o �wHW��f/��o �E��~xv�%��f(�f(�f(��fT5@�f(�f(�f(��%���\U��\]��\���ă��Y��Y��Y��XU��X]��X�f��WX(�(��]��XE��XM��X�f�����f�P�E��D$�G`�X��U��M��$P��������o �E��~@f�E����   �D$�o ��~@�E�Pf�A������$�x �o �E��~h�]�tR�OhW�f/�v(��e�f/�v(�f/�v(��Opf/����v(�f/�v(�f/�v
(���e��\]��\e��\m��U��E�Y��Y��Y��X]��Xe��Xm�f��f�h_^��]� �EW�_^� f�P��]� ���
����U������@�y t�u�u�u�u��U  �E��]� �U�BT��u����\B���^  �y@ �o��   �~��   �D$(u�o��   �~��   �D$(���   W��-P��T$0�|$(�@ �XfW��H(fW��Y�fW�f(��Y��X�f(��Y��X�f/����v
����f(��L$0�X �Y�fW��Y��Y��A8�L$�H�Y\$fW��Y��Y��$�@(fW��X��Y�f(��-���X�f(��\$ �Y��@��\��$�\�(�fT�f(��\��X��Y��Y�f.��L$�T$���Dz�d$�#(�fT��j� �L$W��@��D$f.̟��Dzf(��fT�f(��6� f(�W��\$ f(��X��Y��XL$f.̟��D{1�|$f(��Y,$f(��Y�f(��X��Y��X�f.ԟ��Dz!�E(�����f�@��]� �\�f(�fWP��\��Y��Y��Y��X\$�X��^��^��X��Y��f(ȋEf��f�@��]� ���U���xSVW��� t�u�u�u�uV��R  ��_^[��]� �Mj �X=  �M��j�L=  W�W��M���fE�����E���t8���j S�@@�@8�Ѓ��M���u�uSQ���RH�o �E��~@�E�� ��   ����   ���j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��w`�$���E��%�E���E���E��XE��XE��Yh����W�f/��E�v�M��f/�v(��M������M�� tf(��\�f(��M��W@W��OH�\�f.ȟ��Dzf(���]��\��^�f.ȟ��Dzf(���e��\��^�f.ȟ��Dzf(���u��\��^��GP�� �WX���\�f(�(��Y��gh�Y��Y��X��_`�X��X����Y�f�(��E�f(��Y��YE�(��X��X��X��Gp�D$f��f�`�E�P�����_x��$���w4�o���o)���~a�m�� f�f�@�"%���M����]��E���\���\��\��Y��Y��Y��X��X��X��(�f��(f�`�E��D$���   �$P�����mЃ�,�  �o �~X�E�uf(���M��$ �u�uf(���U��( �e�u(܃8 t W�f/�vf(�f/�vf(�f/�v(؃< t%���f/�vf(�f/�vf(�f/�v(��E��\��\֋E�\��Y��Y��Y����   �X��X�_�X�^�\��\�[�\��Y��Y��Y��X��X��X�f��f�X��]� ������������������U������$  SVW���|$D� t�u�u�u�uV��N  ��_^[��]� �Mj �.9  ��W��L$��u�E� f�@_^[��]� �G@�   �D$0�D$(�\$fD$h;�w1�$�4�   ��   ��_D�É\$%  �yH���@uC�\$�O8fn�������j Q�@@�^ȋ@8�L$h�Ћu��$�   ����uV�t$Q���RH�G8W�f.��o�~P��T$X��$�   ��$�   ��Dz�E�f�P_^[��]� �����$  �^�W���$�   f�$�   f�$�   f�$�   f�$�   ��tjh��$�   VP�� �����  �D$p�C���$�   ��$�   �+��D$H�D$h���ȉ\$���D$8���L$T�D$��I �\$`��fn�����Y��X��D$ ��$�   ���$    �\Ffn�����Y��Y��X���$�   �\N��$�   �\�Y��Y��X��X��ׅ �D$D�H8f/���   �Y�$�   ������j �t$�@@�\ȋ@8�L$(�Ѓ���$�   ��uQ�t$��$�   Q���RH�\$ ��$�   ��$�   ��$�   �Y��Y��Y��XD$8�XL$H�X\$(�XT$0f(���$�   f(��d$8f(��l$Hf(��|$(�t$0�D$ ��D$ �d$8�l$H�t$0�|$(�G�\$`K������D$�V@�L$�\$�L$T�D$�W���W�f/�v ����^��\$X�Y��Y��Y��%�o�$�   �\$X�D$h�l$pf��d$h��$�   �\���$�   �\�����\͋E_�X��X��X�^[f��f�X��]� ������������������U���   VW��� t�u�u�u�uV�J  _��^��]� �uW�f]�W��FT����   �G4���2  �$��#�=���\~�  ����h �]��F���h �]��F���h �Ef]�_�]��}��^f�x��]� �E(��=��_�^f�x��]� �P �o��   �~��   �E��e�u�o��   �~��   �E��e��O4���l  �$�$���   �E��=���H �YM��Y@�X��@(�Y��X�fT@��\��  ��0  ���  �o��  _�~�   �E^�f�x��]� �o�  _�~�   �E^�f�x��]� �8 t&��   ���D$G@$�Q������  ��   �  ��0  ����  �o��   �]��o�(  ��h����o�  �U��o�8  f��Y��o�  �X��E��om�f(���0  �Y��Y��X�(�f��YE��X�f(���   �Y��m���P  �X��X��E��o�H  �8 �YE��M��Ym��Y��X��Y��X��M��oM��U����X�f��X���  ����Y��Y��Y��X��X��X�f(ًEf�_^�f�x��]� ���yn���]�W��U��o@`�o��   ��h����o@p�o��   f��Y��o��   �X��E��om�f(����   �Y��Y��X�(�f��YE��X�f(����   �Y��m����   �X��X��E��o��   ������8 �o�f���   ���(��E��U��Y��Y��Y��X��X��X�f(���������   �@�H �YE��YM��X��@(�Y�3��X�f/�����fn�����$�L������]��}�(�fߋE_^�f�x��]� ��������  q � !D!3#�"� {#����U���@VW��� t�u�u�u�uV�E  _��^��]� �MSj �	0  �M��j��/  W�W��M���fE�����E���t8���j S�@@�@8�Ѓ��M؋�u�uSQ���RH�o �E��~@�E�� [��   ����   ���j V�@@�@8�Ѓ��M؋�u�uVQ���RH�GH��wd�$� &�M��%�M���M���M��XM��XM��Yh�W��M�f/�v
(��M��f/��v����M���M�� t����\�(��M��-���M�f(��E��\��u�f(��e��\ЋE�\�_�\�^�\��\��Y��Y��Y��X��X��X�f��f�h��]� ��%%$%+%U���xVW��� t�u�u�u�uV��C  _��^��]� �u��Sj �'.  j�ΉE�.  j�΋��.  �MW��E�f(��e�Wɋ�fE�����E�fM�fM���tB���j Q�@@�@8�Ѓ��M���u�u�uQ���RH�e�W��o �E��~@�E���t=���j S�@@�@8�Ѓ��M���u�uSQ���RH�o�~`fM�fM��e� [��   ����   ���j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$��*�E��%�E���E���E��XE��XE��Yh�W��E�f/�v
(��E�����f/�v(��E���E����� �e�t�\�(��E�fM؋G4f��u��m��MЃ��  �$��*�  t�M��X���MЃ$ t�U��X���U؃( ��  �}�(��X���  �  tf(��\M���MЃ$ tf(��\U���U؃( ��  f(��\]��  �  t�M��Y���MЃ$ t�U��Y���U؃( �V  �}�(��Y��E  �  W�t)f.���D{�U�f.П��D{
f(��^��f(���MЃ$ t)f.���D{�}�f.����D{
f(��^��f(���U؃( ��   f.����D{�}�f.����D{f(��^��   (��   �  t�M�f/�v
(���MЃ$ t�U�f/�v
(���U؃( tf�E�f/��E�  t�M�f/�v
(���MЃ$ t�U�f/�v
(���U؃( t�E�f/��f���f(��
�U��M��E��\��\֋E�\��Y��Y��Y��G8�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�X��]� d'k'r'y'(V(�(�(�)�)��������U����   S��V�]��{ t�u�u�u�uV�?  ��^[��]� �u��Wj �q)  j�ΉE�e)  �} ������E�W�u�E_^[� f�@��]� �{ ��   ����   ���j W�@@�@8�Ћu�Mă���uVWQ���RH�CH��wd�$��.�M��%�M���M���M��XM��XM��Yh�W��M�f/�v
(��M��f/��v����M���M��{ t����\�(��M���u���W��}j W�@@fE��E�    �E�@8�Ѓ��������uVWQ���RH�K8�Y0��M�o �M��E��~@�E�W���h���f�(���f�8���f�H���f�X�����tjhQ��(���P��y �M����U̍{L�m�3��]�U��m����    �? �  ����̋��������+�fn�����\���Y��X�(�����(���fn�����^��E��E��$�/x �]��,E�j Sfn��������\���YE��X�0�����0����@@�@8�Ѓ���(�����uQS�M�Q���RH�M��M��U��o�]��u���(����~A�M�fօ8����fn�����M��Y��Y��Y��XM��XU��X�(��m��U��]���]�M��M�F����������]��{H tJ��tFfn�W����f.����D{$����^�(��Y��Y��Y�f(�(��f(�(�f(���u��m��e܃{  �K@f(�(��X��m��X��X�uf(Ճ{$ �e�u(܃{( �u�u(��E��\ՋE�\��\�_^�Y�[�Y��Y��X��X��X�f��f�H��]� �+�+�+�+��������U��y Vt�u�u�u�uV��:  ��^]� �Mj �3%  ����t-���j V�I@�I8�у��ȋ�u�uV�uV�RH��^]� �EW�^ �@]� �������������U������(  VW���|$$� t�u�u�u�uV�D:  ��_^��]� �Mj �$  �O@���Y��W��L$�D$�D$�X ��L$0��u�E �@_^��]� ���j Q�@@�@8��W����E���D$xfD$8fD$HfD$XfD$h��tjhP�D$@P�/v ���M����\$@�T$8�t$,��    �T$$���fn�����D$(���YB8�X��D$@fn��BH����YB8�X��D$8�� ��  H��   H�R  9��ta�Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn���M����Y��XD$(��L$��0� ��  �Q�L$<Q�t$�@H��$  Q�����o�~P(�f�f/�vf(�f/�vf(�fn�0��   ��ı t^�Q�L$<Q�t$�@H��$$  Q�����o�~P(�f�f/�vf(�f/�vf(�fn�ı�M����Y��XD$�D$��� �  �Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn������Y��XL$�L$��   ��|� t^�Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn�|��M����Y��XD$�D$���� tL�Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn����+����L$�E���M�T$$��D$(@�D$(���T����t$,�EF�t$,�X������fWP�f(��L$�Y��L$�Y��X��L$0�Y��X��o ����^ȋE_^�\$�D$�d$(f�(��Y\$��$�   ��$�   ����Y��Y��Y��Y��Y��X��X��X�f��f�`��]� �U����y Vt�u�u�u�uV��5  ��^��]� �Mj �   ��W�WɅ�t/���j V�A@�@8�Ѓ��M��u�uVQ���RH�o �~H�E^� f�H��]� U���   VW��� t�u�u�u�uV�;5  _��^��]� �MSj �  ��W���u�E[_^� f�@��]� �uW��M�f�x���fE�fE�fE���tjh��x���VP�cq ��WɃ4�o�~f�E�����e��e��Z  �~T �P  �D& �ȉE�z& j���   P�� ���P��4 �M���o��M�oB�A�M�oB �A �E�oB0�@0�E�oB@�@@�E�oBP�@P�E�Oxf�@fY�@�@(�Y��@(@0���   f�fY�@0�@@�Y��@@@H���   f�fY��YHX@H�HX�E�oG`� �E�~Gpf�@�� ����uP��g���M���o �A`�o@�Ap�o@ ���   �o@0���   �o@@���   �o@P���   �Eƀ�    �Eƀ�    �E�O4���   �E�G@���   �E�GH���   �E�GP���   �E�GX���   �Eǀ�      �Eǀ�       �Eƀ  �8 t
�E���   �< t
�E���   �M̍E�P���   P���   P�uQ�������u�o�x����E��~E�f�E��EP�$ �E����E��   �oP�U��]��\W@�\_Hf.���D{�^��(��oXf.��U���D{�^��(ك8 �]�uYf/�v(��	f/�v(�f/��e�v(��	f/�v(�f/�v(��	f/�v(�f��U��e��8 ��   �< �E���   �����O �]��E������O �]�W�f/�����]�v	�X��]��U�f/�v	�X��U����f/�v�\�(��\��E�f/�vY�\��\��M��J���mO �]��E����`O �U�W�f/�����]�v	�X��U��U�f/�v	�X��U��E�3�9��   �oE�E��E̡����x���Q�E�f�E��@@S�@8�Ѓ���x�����uQS��`���Q���RH[_^�o �~H�E� f�H��]� ���������������U������  ��3ĉ�$�  �ES�]VW���\$(�M�|$ �D$,� t�uPQS����/  �  �HTW�W�f(���  ���  ;GL��  �_@f/���  �H �o��   ��$�   �~��   fք$�   u"�o��   ��$�   �~��   fք$�   �4 W���������,�f�$�  D���$�  f�$  f�$   f�$0  f�$@  f�$P  f�$`  f�$p  f�$�  f�$�  ���   �@0��$�   ��$  (�P��$�  f֌$�  ���   ��P��$�   P��@ �T$8�\$\���o�RTS��$�   �~@��@  �����$  fք$�  fք$�  fք$l  ��$�  Q��$x  ����$�   ��$h  �o��   ��$�   �~��   ��$�   fք$`  fք$H  fք$0  W�fD$p�D$h    f�$�   �D$d    f�$�   Ǆ$�       �$�   fn������$P  ��$8  ��$   �@�$QR��   ��$�   Q�Ѓ��o�~@�D$P�\$(�D$HfL$0���  ����\$,�@	��   ��$�   �|$P��$�   ��$   �ST����Y�W�Yˍ�@  Q�YӍ�$�   ���\$p�X��D$x�X���$�   �X�f�fn������$�   f֌$�   ��$P  f֌$`  ��$8  f֌$H  ��$   f֌$0  �@�$QR��   ��$�   Q��������o�~@�D$PfL$0��������|$ �\$(�D$H�G4H��   H�H  9D$T�8  �T$`�D$h�\�$�   �\�$�   �L$p�\�$�   �Y��Y��Y��X��X��e ���D$G8$�B����荄$�   �OP����\$(�D$(�$P��� ���@�$�q�|$T ��   �T$`�D$h�\�$�   �\�$�   �L$p�\�$�   �Y��Y��Y��X��X��|d ���D$G8$����������$�'���D$8���\$ �L$ f�fY�D$0�D$H�Y�fL$0�W�W��f�C��$�  ��_^[3��I ��]� ��������������U���|S��V�]��{ t�u�u�u�uV�*  ��^[��]� W�}W�fE��E�OT����  �{@ �o��   �E��~��   f�E�u�o��   �E��~��   f�Eġ��Q�@�@X��3ɉE���M����  ���Q�wT�@�@T�Ѓ����{L �u�t8������   �M�RT���v�KLP� 3�9SH��3Ƀ����;��   �GT���   ��@  ���}��]����   �]���   ���   ����{T�]��@��(  �}���p  W�}jSRQ�M�Q�OTV�u�Q�M�Q�Ћ]���,�o �{D �~X�E��C8�M��U��Y��Y��Y��X]��XM��XU�th���f(�W��e�f/�v�]��f/�v�E�f/�v(��	f/�v(�f/�v(�f��M��#f/�v(�f��M���M��U��]�MA�M;M��y����E�oE�_^� [�E�f�@��]� ����U���0VW��� t�u�u�u�uV�>(  _��^��]� �Mj �  ����u�EW�_^ �@��]� ���j V�@@�@8�Ѓ��M��u�uVQ���RH�oE�G4�M�W�����EЃ�w&�$��B�E��E���M���]���U�G8�E��eЃ�w(�$��B�e���E���M���]���U��G<��w�$�C(��(��(��(ʋE�oE�_^� f�H��]� �_B@BLB_BSBZBxBB�B�B�B�B�B�B�B�B�B�B����U����   SVW���}�� t�u�u�u�uV�&  ��_^[��]� �]W�W��{T �	  �Mj ��  (�������U�f�4�����t=���j V�A@�@8�Ѓ��������uSVQ���RH�o ��4����~@�E��P W��KTW�fE��M��o��   �E��~��   f�E�u�o��   �E��~��   f�E��G@3�9��  �Y`���3�9WTQD�3��E��X�����u�@�E��@X�Ѓ�����  �E��E��E��E���I ���V�sT�@�@T�Ћ؃��]؃�$   �n  �\ t8������   �M�@T���s�O\P� 3�9WX��3Ƀ����;��0  �GH�]�U��M��e��[T�Y�j �Yȍ�@  ������   ���   �Y����   j���   �X��X�W��X��   �M��]��E�W�f�|����e�f�d�����t�����(  ���   �@��V�u��u؋�d  WRQ�M�Q�M�Q��d���Q��|���QVS�Ѓ�8���S  �}���  �E�    �E�    �9 t$�E�P�E�P�GT��0  Q�? ���}� �  ���   ��   ���W��WTW�f����f�L����E���,�����\����H��L���P�����P��(  ���   P�E�P�E�P���   ��P��`  ���$j jVR����L�����4��T�����\����Y�|����}��YU��Y]��G8�Y��Y��Y��XM��XU��X]��M��U��]��,  ��l�����d���f(��M�f(��e���t����U��Y��GT�Y܋��   �X�f(��Y��X��@ �Y���Y��Y��Y��\��H�\��\��Y��Y��X��H(�Y��X�W�f/���   �M��nN f(�W�f(�f(��YM��Y�|����YU�f/�vf(�f/�vf(�f/�vf(؋}��G8�Y��Y��Y��E��X��E��E��X��E��E��X��E���}�����]�E�@�sT�@X�Ћu��;��H����E��M��
�M��E��Y�4����Y�<���f(��E��YE�fыE_^[�f�@��]� �����������U��y Vt�u�u�u�uV�T!  ��^]� �q4�M�  ����u�EW�^ �@]� ���j V�@@�@8�Ѓ��ȋ�u�uV�uV�RH��^]� �������������U����y t�u�u�u�u��   �E��]� �I4��t1����U��uR�@ �@X�ЋM�o ��~@��f�A��]� �EW� �@��]� ��������������U����   �y Vt�u�u�u�uV�N   ��^��]� �u��SWj �
  j�΋��
  j�΋��
  j�ΉE�
  �uW��E�W��M�fE�fE�fE�fE���tjh��|���VP�m\ ����E��E����1> �Fݝ|����E��E����> �%��W�f/��|����]�v�X�f/F�U�v�X����3�3�f/ٍQrf/�G�f/�rf/�GA���m  �$�@L���^  ����E��Y�W�Y��Y���|����U��E��"������|����uQW��d�����   ���  ����E��Y�S�Y��Y��\��U��E���|�����!������|����uQ������   �]����   ����E��Y�S�Y��Y��\���|����E��U��j!������|����uQ��4����S�]��tc����E��Y�S�Y��Y��\��\��E���|����U��!������|����uQ��L���S�Q���RH�o fE��~@�EfM�_[�^f�@��]� ��JKfK�KU���   VW��� t�u�u�u�uV�  _��^��]� �G`W����f.����Dz�W`�Ghf.����Dz�Wh�Mj �  ����u�EW�_^ �@��]� �EW��G8�%P�f.��o��U��]��\Wp�\_x�U��]���D{	fW��U��G@f.����D{	fW��]��GX�.T �E��GX�D �oe���`���f(��E�f(�f(��YU�jh�YE��Y��Y��\��X��^_`�^Wh�\_H�XWP�X_p�XWx�}WP�]��U���X �oM����E�f��~G��`���j fօp����@@V�@8�Ѓ���`�����uQV�u��V�RH_��^��]� ���������������U��y t�u�u�u�u��  �E]� �EW� �@]� �������������U��E�A�E    ]�*�  ����������U����SV�u�ً@@WV�@,�Ћ�����΋����   �RT�ҋ��j Ph�  �Q�ϋBl�Ћ����j h�  �Q�ϋ��   �ҋ���u
_�s^[]� ����΋��   �@��=�� u
_�s^[]� ����΋��   �@��=�� t����΋��   �@��=�� u���  P蚷������P�  �C_^[]� �����U��W�f/Ev����E�E]�����E�E]��������������������������������U���X����M�SVQ�@�@�С���M�j j�hp��@Q�@�С���M�E�    ���@�@<�Ћ���؍E�P�I�I�ы��j j�h���A�M�Q�@�С���M����@j�Q�M�@DQ�M�Ћ�����E�P�I�I�у�����  W�}��C�;�u}����M�Wj Q�@�M�@P�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���MQ�M�Q�@�@�С���M�Q�@�@�Ѓ��-  G;��$  ��$    ����M�jWQ�@�M�@P�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M����E�    �@j Q�M�@@Q�M��Ѕ�����@��   �u��@P�M�j Q�M�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���MQ�M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@��G�� ;��������@�M�Q�Ѓ�_����uV�@�@�С���MVQ�@�@�С���H�E�P�I�ы���EP�I�I�у���^[��]� ���������������V���hS  �t��ݏ  j jjZjZ�ȉF0諌  �N0j j j 荍  �F    ���F   �F    �F   �F   �F    �F    �F$   �F(   �F,    ^����VW��j j h,� �t��^ �O0�w0���j�  V�T�  ����_^��R  ��������U����SV���   �@(�Ћ]����t\W��tT���V�@@�@,�Ћ���������   �΋RT�ҋ��h*� Ph�� �Q�ϋBl��;�tj ����������u�3�_^[]� _��^[]� �������U����SV���   �@,�Ћ]����t\W��tT���V�@@�@,�Ћ���������   �΋RT�ҋ��h*� Ph�� �Q�ϋBl��;�tj ����������u�3�_^[]� _��^[]� �������U����V��W�@@V�@,�Ћ�����΋����   �RT�ҋ��j PkEd�Q���� P�Bl��_^]� ������   �@x��U��} �   V�   E���Q�@@�@��#�3Ƀ�;�����^]� ���������̡��V��V�@@�@�Ѓ��u���V�@@�@�Ѓ��u3�^ø   ^��������̡��V��W�@@V�@,�Ћ�����΋����   �RT�ҋ��h*� Ph�� �Q�ϋBl��_^���������U���0���Q�@@�@,�Ћ����W���fE��E��A�M�Qh�� �MЋ��   Q�����o�~@�Ef�E���Ef����]� ����U���0���Q�@@�@,�Ћ����W���fE��E��A�M�Qh�� �MЋ��   Q�����o�~@�Ef�E��f��H��]� �����̡��Q�@@�@,�Ћ�����ЋA��j h=  ���   �����U������ �@@VWQ�@,�Ћ�����E�P�I�I�ы�����A�M�Qh;  �M����   Q���Ћ�����}W�I�I�ы��WV�A�@�С���H�E�P�I�ы���E�P�I�I�у���_^��]� ���������������U������ �@@VWQ�@,�Ћ�����E�P�I�I�ы�����A�M�Qh<  �M����   Q���Ћ�����}W�I�I�ы��WV�A�@�С���H�E�P�I�ы���E�P�I�I�у���_^��]� ��������������̡��Q�@@�@,�Ћ�����ЋA��j h>  ���   �����U������ �@@VWQ�@,�Ћ�����E�P�I�I�ы�����A�M�Qh?  �M����   Q���Ћ�����}W�I�I�ы��WV�A�@�С���H�E�P�I�ы���E�P�I�I�у���_^��]� ��������������̡��V�񋀈   �@T��j P���y  ^��U����VW���@@W�@,�Ћ����kMd���B�u���� Q�@p���Ѓ} tjW���  j j h,� �zX ��_^]� �U�������   �@|]��������������U��} �   SVW�   ��E�����} Stw�@@�@��#ǃ�;�t���S�p@�F���P�FS�Ѓ��} t\����ˋ��   �@P�Ћ���tD������   �ˋRL�ҋ��S���   �΋@h��_^[]� �p@�F����#�P�FS�Ѓ�_^[]� �������U����Q�@@�@,�Ћ�����ЋA���uh�� �@p��]� ��������������U������Q�@@�@,���E��������E��E�E�W��E��A�M�Qh�� �ʋ@H�Ћ�]� ������������U������Q�@@�@,��E�������E�W��E��A�M�Qh�� �ʋ@H�Ћ�]� ��������U����V��V�@@�@,�Ћ�����ȋB�uh=  �@0��jV���w  j j h,� �YV ��^]� �U����Q�@@�@,�Ћ�����ЋA���uh;  �@8��]� ��������������U����W��W�@@�@,�Ћ�����ȋB�uh>  �@0�Ѓ} t
j W����  j j h,� ��U ��_]� �����������U����Q�@@�@,�Ћ�����ЋA���uh?  �@8��]� �������������̡��VW���@@W�@,�Ћ�������΋Rj h=  ���   �ҋ���Q3Ʌ����B0Qh=  ����jW���(  j j h,� �
U ��_^����̡��SV�ً@@WS�@,�Ћ�������ϋRj h>  ���   �ҋ�����Q3Ʌ����R0Qh>  ���҅�u	VS���   j j h,� �T ��_^[��������������U����Q�@@�@�ЋЃ�#U3�;U��]� �����������U����VW���p@W�F��EP�FW�Ѓ�_^]� ��������U����VW���p@W�F�ЋU��#�P�FW�Ѓ�_^]� ����U������4�@SV�ٍM̋@WQ�С���$��u��j j��H��D�P�E�P�A�С���M�Q�@�@�С���M�j j�h,��@Q�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M��4�@�@<�Ћ��j�j��Q�M�QP�M�BL�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С���}W�@@�@,�Ћ�����ЋA��jh�  �@0�С���ϋ��   �@��-�� �Q  ���@  ��&�7  ���7  ����ϋ��   �@P�Ћ���Ћ��   �ʋ@X�Ћ؅��  ��    ���j S�A@�@8�Ћȃ�3��M��E��� �P�R\��tZ���S�@@�@,�Ћ���������   �ˋRT�ҋ��j PV�Q�ϋBl�Ћ};�u�����j hȴ ���   �@�ЋE��d�M�@�E��Q� |����W�@@�@,�Ћ���������   �ϋRT�ҋ��h*� Ph�� �Q�΋Bl��P��������؅�����_^[��]� W���   _^[��]� �������U��V�gE ������u�I@�I,�у���Vh�  ��l  �Ѕ���   ������   �ʋ��   �Ћ�����   W���$    ����΋��   �@��=.� ug���V�@@�@,�Ћ�������Q��j h�  ���   �ҋ���P3���?B OЋARh�  �ϋ@4�С����j j���   �@�С���΋��   �@(�Ћ����d���_^]� ��������������U������V�uV�@@�@,�Ћ��W����E���fE�A�M�Qh�� �ʋ@H�С��V�@@�@,�Ћ�������Q��j h�  �R0�ҋ��jh�  �A�΋@0�С����j h�  �@�@4�С����jh5  �@�@0�С����jh6  �@�@0�С����jh7  �@�@0�С����j h8  �@�@0�С����j h:  �@�@0�С����jh9  �@�@4�С���M�Q�@�@�С���M�j j�hx��@Q�@�С���M����@Qh;  �΋@8�С���M�Q�@�@�С�����΋@j h=  �@0�и   ^��]� ������U��]�Gs  �������U��]��s  �������U��Q���S�u�M��@@�@,�ЋM����j �9� ���������w �����j h8  �@���   ��[��]� �u�M��u�u�u�u�us  [��]� ��������������U������SVW�@@�ً}j W�@8�Ћu���E���(  t��tA���M  ���D  �����j hȴ ���   �@��j j h,� �M ���  �M�	�; ����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�ЋE���Wj*�; ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�ЋE����; ����M�Q�@�@�С���M�j j�h��@Q�@�С���M�Q�@�@�Ѓ��5��-�� t��u'jW�����������ϋ��   �@T�ЋMP��Rh�u��VW�Gq  _^[��]� ��������������U������S�]V���   �M���W�@�Ћ}=�� �����   ���   �ϋ@T�Ћ��(@ ;�ug����M�Q�@�@�С���M�j j�h���@Q�@�С���M�Q�@�@�Ћu�����j W����������j h�� ���   �@����u��u���uWS�u�xp  _^[��]� �@@W�@,�Ћ�����؋��   �ϋ��   �ҋЅ�tH����uj ���   �ʋ �Ћ����j V�ϋ��   ���   �ҋ��Vh�  �A�ˋ@p��_^�   [��]� ���������������U��Q���SVW�@@�}j W�@8�Ѓ��E�3۾�� ���S�R\��tj���W�@@�@,�Ћ���������   �M�RT�ҋ��j PV�Q�ϋBl�Ћ���t&���j W�I@�I8�у��ȋ�u�uW�RD��u�}��dC��Q� }�E��v���3�_^[��]� ����U��Q���SVW�@@�}j W�@8�Ѓ��E�3۾�� ���S�R\��t`���W�@@�@,�Ћ���������   �M�RT�ҋ��j PV�Q�ϋBl�Ћ���t���j W�I@�I8�у��ȋW�RL�}�E���dC��Q� |�_^[��]� �����U��V�u�u���uV�{������u  ���SWj �@@V�@8�Ћ����V�I@�I,�ы�������Q��j h�  ���   �҅��'  �����jh�  �@�@0�С����j h=  �@���   �ЉC�ϡ��jh�  �@���   �ЉC�ϡ��j h�  �@���   �ЉC�ϡ��jh9  �@���   �ЉC�ϡ��jh8  �@���   �ЉC�ϡ��j h:  �@���   �ЉC�ϡ��jh5  �@���   �ЉC �ϡ��jh6  �@���   �ЉC$�ϡ��jh7  �@���   �ЉC(������   �@T���ЉC,_3�[^]� ���������U����VW�}�@@j W�@8�Ѓ��ȋ�Rd��~r���W�@@�@,�Ћ�����ϋ����   �RT�ҋ��j Ph�� �Q�΋Bl�Ћ���t.���j V�I@�I8�у��ȋ�u�uV�uV�RH_��^]� �EW�_^ �@]� ����U��V�u��V��������V�@@�@,�Ћ�������Q��j h�  ���   �҅�t�����j h�  �@�@0��^]� �����U���@V�  (���M����E�fE�P� ��E��,������M�Q���   �@@�Ћ�����Q��Ph�  �E�P���   �Ћ���u�o ���   ��~@�E��	Pf�F�у���^��]� ���̸   �����������U����V�uV�@�@�Ѓ}c���j j��I�Iuh��V�у���^]� h$�V�у���^]� ̸   � ��������U��MW��E�A��c��   ���l�$��l(�����p��f�I]� (`�������f�I]� (P�������f�I]� (p��0��f�I��]� �Klil�l�l�l ����3���������������U����   SVW�}���u�8 ���^�]����  �N0����  ���Q�@�@�Ѓ�����  ���k������q  ���S�@@�@,�Ћ�����؋Q��j h�  ���   �҅��<  �����j h�  �@�@0�ЋN0�p  �N0j jjZjZ�Pq  �N0j j j �2r  W������WfE��E��  ������jQ�u���PD����  ������  �@�W��E�3��E�    f�E�fE��E�   ��x�������]�f�E��fn�3�����^��M����$    �d$ fnÍ�`�������jQ�M��u�^�Q��f���`���W�fօp����PH���W��of/�f]��~Pv�M��f/�v�E���]��]�f/�v�M��f/�v�E���]�f/�v(��	f/�v(��oE����M�f�U��E�j�@Q�M�Q���  ���p��ofM��~@����E��YH�,�(�f�P�Y��Y��,�P�,�P��  WS�v0���M�C�@���$��Z�����G��Z���������u�PL��$����9  _^[��]� ���������U����j �u�@@�@8�Ѓ�]�������U��E���   ����V��i�|  ��Hs�$��r�E^�    �@   ��]ËE^�    �@   ��]ËE^�    �@   ��]ËE^�    �@�   ��]ËE^�    �@    ��]ËE^�    �@x   ��]ËE^�    �@   ��]ËE^�    �@
   ��]ËE^�    �@    ��]�(���EЋMfE�P����E��&���E^��]�(`���p����Mf�p���P����E���%���E^��]�(��E��MfE�PW��E��%���E^��]�(p���@����Mf�@���P�����P����t%���E^��]�(���E�MfE�P����E��G%���E^��]�( ��E��MfE�P�(��E��%���E^��]�(0��E��MfE�P����E���$���E^��]�(����X����Mf�X���P� ���h����$���E^��]�(����(����Mf�(���P�H���8����$���E^��]ËE^�     �@    ��]�yp�p�p�p�p�p�pqcq�q!q6q�q�q!rNr{r�r�r  	
��������������U���\V�? �����h&� �A�ʋ@T�Ћ�����  �M��X  ���t? �����Vh&� �A�ʋ@D�ЍM���X  �O? �����h&� �A�ʋ@T�Ћ���u^��]á���M��E�   �E�   Q���   �@8�Ћ�����Q��PhM  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��PhR  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��RhN  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����QP�B4��hO  �С���M�Q���   � �С���M��E�   �E��   Q���   �@8�Ћ�����Q��PhP  �B4�С���M�Q���   � �С���M��E�   �E�    Q���   �@8�Ћ�����Q��PhQ  �B4�С���M�Q���   � �С���M��E�   �E�x   Q���   �@8�Ћ�����Q��PhS  �B4�С���M�Q���   � �С���M��E�   �E�   ���   �@8Q�Ћ������ҋA��Rh]  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��PhT  �B4�С���M�Q���   � �С���M��E�   �E�
   Q���   �@8�Ћ�����Q��PhU  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��Rh\  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��Ph_  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��RhZ  �΋@0�С���M�Q���   � �С���M��E�   �E�    Q���   �@8�Ћ������ҋA��Rh[  �΋@0�С���M�Q���   � �Ѓ�(���E�fE��M����P�E��������M�Q���   �@@�Ћ�����Q��Ph^  �BH�С���M�Q���   � ��(`��E����M�fE����P�E��+������M�Q���   �@@�Ћ�����Q��PhW  �BH�С���M�Q���   � ��(��E����M�fE�W�P�E���������M�Q���   �@@�Ћ�����Q��PhX  �BH�С�����   �M�Q� �С���M��E�   �E�   Q���   �@8�Ѓ��M�fn�������QhY  ��f�E��E��@�@H�С���M�Q���   � ��(p��E����M�fE����P�E���������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE����P�E��������M�Q���   �@@�Ћ�����QP�BH��h�  �С���M�Q���   � ��( ��E����M�fE��(�P�E��+������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(0��E����M�fE����P�E���������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE�� �P�E��[������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE��H�P�E���������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � �Ѓ���^��]����������U�����MQ�@�@�Ѓ�]��������U��V��W��F�N����F�-+  �u����  ��^]� ������������U��VW��j j h,� �t��4 �O0�w0���Wa  V�Ae  �����(  �Et	W�[!  ����_^]� U����Af.���E����Dz���]���u���]���̡�����   �@(�������   �@,�������   �@x����Q�@@�@�����������������U���0���Q�@@�@,�Ћ����W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�Ef�E���Ef����]� ����U���0���Q�@@�@,�Ћ����W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�Ef�E��f��H��]� �����̡��Q�@@�@,�Ћ�������Q�$�A��h�  ���   ������������U���0���Q�@@�@,�Ћ����W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�E�,�fɉ�E�,�f�E����]� U���0���Q�@@�@,�Ћ����W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�Ef�E��f��H��]� ������U����Q�@@�@,�Ћ���Ѓ��A�Mj ���   �����  ��Q����]� �U�������   �@|]��������������U����VW���p@W�F�Ѓ} t������P�FW�Ѓ�j j h�� �U1 ��_^]� ������������U������Q�@@�@,��fnE�����������E�fnE����E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ����U������Q�@@�@,��E�������E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ��������U����Q�@@�@,�Ћ�����EQ�$�A��h�  �@,��]� ���������U������Q�@@�@,��fnE�����������E�fnE����E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ����U������Q�@@�@,��E�������E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ��������U������VWQ�@@�@,�Ћ�����u���A�Nd�����@0j Q���С���4�W���fE��E��P�E�P���  P�BH�С��������ϋP���  �$P�B,��_^��]� ������������U������P�@@VWQ�@,�Ћ�����u���A�Nd�������   j Q���Ѕ���   ����4�W���fE��E��P�E�P���  P�E�P���   �Ѓ����o �E��~@���f�E�����$�P���  P���   �С�����]��E��ϋ@�$h�  �@,�С���M�Qh�  �ϋ@�@H��_^��]� ��������U���P���VWQ�@@�@,�Ћ����W���fE��E��A�M�Qh�  �M����   Q���Ѓ����o �E��~@���f�E�����$�@h�  ���   �С���ϋuj�]��P�Fd����P�B0�С���4��ϋP�E�P���  P�BH�С�����E��ϋP���  �$P�B,��_^��]� ��̸   � ��������� �������������U��E���   ����V��i�|  ����$����E^�    �@   ��]ËE^�    �@   ��]ËE^�    �@   ��]ËE^�    �@�   ��]ËE^�    �@    ��]ËE^�    �@x   ��]ËE^�    �@   ��]ËE^�    �@
   ��]ËE^�    �@    ��]�(���EЋMfE�P����E��e���E^��]�(`���p����Mf�p���P����E��2���E^��]�(��E��MfE�PW��E��
���E^��]�(p���@����Mf�@���P�����P��������E^��]�(���E�MfE�P����E�����E^��]�( ��E��MfE�P�(��E��z���E^��]�(0��E��MfE�P����E��M���E^��]�(����X����Mf�X���P� ���h�������E^��]�(����(����Mf�(���P�H���8��������E^��]ËE^�     �@    ��]��.�C�X�m��������6���օ^�������Q���  	
��������������U���\V�+ �����h&� �A�ʋ@T�Ћ�����  �M��D  ����* �����Vh&� �A�ʋ@D�ЍM��DD  �* �����h&� �A�ʋ@T�Ћ���u^��]á���M��E�   �E�   Q���   �@8�Ћ�����Q��PhM  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��PhR  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��RhN  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����QP�B4��hO  �С���M�Q���   � �С���M��E�   �E��   Q���   �@8�Ћ�����Q��PhP  �B4�С���M�Q���   � �С���M��E�   �E�    Q���   �@8�Ћ�����Q��PhQ  �B4�С���M�Q���   � �С���M��E�   �E�x   Q���   �@8�Ћ�����Q��PhS  �B4�С���M�Q���   � �С���M��E�   �E�   ���   �@8Q�Ћ������ҋA��Rh]  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��PhT  �B4�С���M�Q���   � �С���M��E�   �E�
   Q���   �@8�Ћ�����Q��PhU  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��Rh\  �΋@0�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ�����Q��Ph_  �B4�С���M�Q���   � �С���M��E�   �E�   Q���   �@8�Ћ������ҋA��RhZ  �΋@0�С���M�Q���   � �С���M��E�   �E�    Q���   �@8�Ћ������ҋA��Rh[  �΋@0�С���M�Q���   � �Ѓ�(���E�fE��M����P�E���	������M�Q���   �@@�Ћ�����Q��Ph^  �BH�С���M�Q���   � ��(`��E����M�fE����P�E��	������M�Q���   �@@�Ћ�����Q��PhW  �BH�С���M�Q���   � ��(��E����M�fE�W�P�E��(	������M�Q���   �@@�Ћ�����Q��PhX  �BH�С�����   �M�Q� �С���M��E�   �E�   Q���   �@8�Ѓ��M�fn�������QhY  ��f�E��E��@�@H�С���M�Q���   � ��(p��E����M�fE����P�E��[������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE����P�E���������M�Q���   �@@�Ћ�����QP�BH��h�  �С���M�Q���   � ��( ��E����M�fE��(�P�E��������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(0��E����M�fE����P�E��#������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE�� �P�E��������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � ��(���E����M�fE��H�P�E��S������M�Q���   �@@�Ћ�����Q��Ph�  �BH�С���M�Q���   � �Ѓ���^��]����������U����M�������E���u��]� SV�u��Wj �6� j �΋��+� �u��؍E�V�u�7P�G����M���P�3�i� ����M�Q���   � �Ѓ��   _^[��]� �����U���V��M�hM  �ڂ ��M�j Q���PD�M��Մ hR  �M�踂 ��M�j Q���PD�M�賄 hN  �M�薂 ��M�j Q���PD�M�葄 hO  �M��t� ��M�j Q���PD�M��o� hP  �M��R� ��M�j Q���PD�M��M� hQ  �M��0� ��M�j Q���PD�M��+� hS  �M��� ��M�j Q���PD�M��	� h]  �M��� ��M�j Q���PD�M��� hT  �M��ʁ ��M�j Q���PD�M��Ń hU  �M�訁 ��M�j Q���PD�M�裃 h\  �M�膁 ��M�j Q���PD�M�聃 h_  �M��d� ��M�j Q���PD�M��_� hZ  �M��B� ��M�j Q���PD�M��=� h[  �M�� � ��M�j Q���PD�M��� h^  �M���� �j �M�Q���PD�M���� hW  �M��܀ ��M�j Q���PD�M��ׂ hX  �M�躀 ��M�j Q���PD�M�赂 hY  �M�蘀 ��M�j Q���PD�M�蓂 h�  �M��v� ��M�j Q���PD�M��q� h�  �M��T� ��M�j Q���PD�M��O� h�  �M��2� ��M�j Q���PD�M��-� h�  �M��� ��M�j Q���PD�M��� h�  �M��� ��M�j Q���PD�M��� h�  �M��� ��M�j Q���PD�M��ǁ �   ^��]� �����������U������S�M��M�W�@Q�@�С���M�j j�h,��@Q�@�Ћ}�E����P�Y� ���M���Q�Ë@�@�Ѓ���t
_3�[��]� V�u� �  hM  �M�� �]��M�WQ�ˋ�PD�M��� hR  �M���~ ��M�WQ���PD�M���� hN  �M���~ ��M�WQ���PD�M��π hO  �M��~ ��M�WQ���PD�M�讀 hP  �M��~ ��M�WQ���PD�M�荀 hQ  �M��p~ ��M�WQ���PD�M��l� hS  �M��O~ ��M�WQ���PD�M��K� h]  �M��.~ ��M�WQ���PD�M��*� hT  �M��~ ��M�WQ���PD�M��	� hU  �M���} ��M�WQ���PD�M��� h\  �M���} ��M�WQ���PD�M��� h_  �M��} ��M�WQ���PD�M�� hZ  �M��} ��M�WQ���PD�M�� h[  �M��h} ��M�WQ���PD�M��d h^  �M��G} ��M�WQ���PD�M��C hW  �M��&} ��M�WQ���PD�M��" hX  �M��} ��M�WQ���PD�M�� hY  �M���| ��M�WQ���PD�M���~ h�  �M���| ��M�WQ���PD�M��~ h�  �M��| ��M�WQ���PD�M��~ h�  �M��| ��M�WQ���PD�M��}~ h�  �M��`| ��M�WQ���PD�M��\~ h�  �M��?| ��M�WQ���PD�M��;~ h�  �M��| ��M�WQ���PD�M��~ ��]����VW�u�F>  ^_[��]� �������������U���   SVW���]����}�؅��/  j ���~ ���������i�  ��l��$�\�j ���~ �0�E�P�������P���   �@8�Ѓ��ϋ�j �T~ ���V�0�Q�ˋ��   �ЉE�M����E�   j Q���   �u�@�С���M�Q���   � �ЍM����Q���   � �ЋE����   _^[��]� j ����} �0�E�P����������p���j �ϋ��} ���V�0�Q�ˋ��   �ЉE؍MС���E�   j Q���   �u�@�С���M�Q���   � �ЍM��\���j ���X} �0�E�P�}������P���   �@@�Ѓ��ϋ�j �-} ���V�0�Q��p���P�ˋ��   �ЍM�Q�M��o Q�E��~@���f�E��E�    �E�    ���   �@�С���M�j Q�u���   �@�С���M�Q���   � �С���M�Q���   � �ЋE����   _^[��]� �u���uW�u��;  _^[��]� �I 8��_�?�          ����������U��SVW���s����}�؅���  j ���{ ���������i�~  ��ȝ�$�������u���   �@8�Ѓ��ϋ�j �}{ ���V�0�Q�ˋB4�ЋE_^[��   ]� ����u���   �@8�Ѓ��ϋ�j �7{ ���V�0�Q�ˋB0�ЋE_^[��   ]� �M�����j �ϋ���z ���V�0�Q�B0����j j h,� �E��� ���   _^[]� ����u���   �@8�Ѓ��ϋ�j �z ���V�0�Q�B4맡���u���   �@@�Ѓ��ϋ�j �vz ���V�0�Q�BH�r����M����j �ϋ��Oz ���V�0�Q�ˋBH��j j h˴ �K����u���uW�u�9  _^[]� ��"�h���)���^���  ��������������U�����E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW� ������u_^]�Wj V�F ��������F�H�   _^]�������������U��M��t+�=H� t�y���A�u	�E]�� ����@�M� ]��]����������U��M��t+�=H� t�y���A�u	�E]� ����@�M� ]��]����������U�����E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW� ������u_^]�Wj V�F ��������F�H�   _^]�������������U�����E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW� ������u_^]�Wj V�� ��������F�H�   _^]�������������U�����E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW� ������u_^]�Wj V�F ��������F�H�   _^]�������������U�����u�@� �Ѓ�]����������U�����u�@� �Ѓ�]����������U��M��t����@�M��@  ]��]á��hﾭދ@��@  ��Y����������U��V�u���t���Q�@� �Ѓ��    ^]�����������U�����@���  ]��������������U��E��t�x��u�   ]�3�]������U�����@��  ]�������������̡���@��   ��U�����E��t!�u�I�   �u;�B�P���   �Ѓ�]ù   ;�VB�W�xW�� ������u_^]�Wj V�
 ��������F�H�   _^]�����������U��M�   �����Dʅ�t�u�@�uQ���   �Ѓ�]Ã�VB�W�yW�s ������u_^]�Wj V�)
 ��������F�H�   _^]����������������U�����u�@� �Ѓ�]����������U�����u�@� �Ѓ�]����������U��E�   ;�VB�W�xW�� ������u_^]Ã} tWj V�	 ��_������F�H�   ^]����������������U�����E��t;�} �   �u�I�ut;�B�P���   �Ѓ�]Ã�B�P���  �Ѓ�]ù   ;�VB�W�xW�4 ������u_^]Ã} tWj V�� ��_������F�H�   ^]�����������U��M�   �����Dʅ�t*�} �u�@�uQt���   �Ѓ�]Ë��  �Ѓ�]Ã�VB�W�yW� ������u_^]�Wj V�V ��������F�H�   _^]�������������U�����u�@� �Ѓ�]����������U�����u�@� �Ѓ�]����������U����Q���   �@X�Ћȃ���u]� ����u�u�@|Q�@�Ѓ�]� ����U����Q���   �@X�Ћȃ���u]� ����u�u�@|Q�@8�Ѓ�]� ����U��UV��j j j ����R�@�@�Ѓ��F��^]� ���̡��Vj ��@j j �6�@�Ѓ��F^�U��V��N��u3�^]� ���Q�u�@�u�6�@�Ѓ��F�   ^]� �������������������������������̅�t�j������̡���@��  �����@��(  ��U�����U���@R��   �ЋMP�m  �M��  �E��]� �����������̡���@��$  ��U�����@��  ]��������������U�����@���  ]�������������̡���@��  ��U�����@���  ]��������������U�����@��x  ]��������������U�����@��|  ]�������������̡���@��d  ��U�����@��p  ]��������������U�����@��t  ]��������������U���EV�����t	V��������^]� �������������̡���@$�@X�����U�����@$�@\]�����������������U�����u�u�@$�uQ�@`�Ѓ�]� ��������������̡��V��V�@�@�С��V�@$�@D�Ѓ���^�����������U����V��V�@�@�С��V�@$�@D�С���uV�@$�@d�Ѓ���^]� ���U����V��V�@�@�С��V�@$�@D�С���uV�@$�@�Ѓ���^]� ���U����V��V�@�@�С��V�@$�@D�С��V�u�@$�@L�Ѓ���^]� ��̡��V��V�@$�@H�С��V�@�@�Ѓ�^�������������U�����uQ�@$�@L�Ѓ�]� �����U�����@$�@]����������������̡��Q�@$�@�Ѓ����������������U�������@$VWQ�@�M�Q�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]� ���U�����uQ�@$�@�Ѓ�]� �����U�������@$VWQ�@ �M�Q�Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у� ��_^��]� ����U�������@$VWQ�@$�M�Q�Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у� ��_^��]� ����U���,�E�VWP�o������P�E�P�I$�A�Ћ�����}W�I�I�ы��WV�A�@�С���M�Q�@�@�С���H$�E�P�IH�ы���E�P�I�I�у� ��_^��]� ������̡��Q�@$�@(��Yá��Q�@$�@h��Y�U�����uQ�@$�@,�Ѓ�]� �����U�����uQ�@$�@0�Ѓ�]� �����U�����uQ�@$�@4�Ѓ�]� �����U�����uQ�@$�@8�Ѓ�]� �����U�����u�u�@$Q�@P�Ѓ�]� ��U�����uQ�@$�@T�Ѓ�]� �����U�����@$�@l]����������������̡���@$�@p�����U����V��V�@$�u�@L�Ѓ���^]� ���������������U����V�uV�@�@�С��V�@$�@D�С��V�u�@$�@L�Ћ���uV�I$�I@�у���^]���U����V�u��@$V�@@�Ѓ���^]� ���������������U�����uQ�@$�@<�Ѓ�]� �����U�����uQ�@$�@<�Ѓ����@]� U�����@(�@]����������������̡���@(�@�����U�����@(�@]�����������������U�����@(�@]�����������������U�����@(�@ ]�����������������U����j�u�@(�u�@��]� ����U�����u�u�@(�u�@$��]� ��̡���@(�@(����̡���@(�@,����̡���@(�@0�����U�����@(�@4]�����������������U�����@(�@X]�����������������U�����@(�@\]�����������������U�����@(�@`]�����������������U�����@(�@d]�����������������U�����@(�@h]�����������������U�����@(�@l]�����������������U�����@(�@p]�����������������U�����@(�@t]�����������������U�����@(�@x]�����������������U�����@(���   ]��������������U�������@V��M�Q�@�Ѓ��E���P�   ��u3������M�Q�u�@$�@�Ѓ��   ����E�P�I�I�у���^��]� ������U��Q����U�R�@(�@X�Ѕ�u��]� �E3�8M�����   ��]� ���������U�������E�    �E�    V�@(��M�Q�΋@h�Ѕ�t�M������u@�@�M�Q�@�С���M��uQ�@�@�С���M�Q�@�@�Ѓ��   ^��]� �@h��he  Q���   �Ћȃ�����M��@(��u�@4��j���3�^��]� �@j �u�Q���Ѕ�u�E�P������3�^��]� ���j �H�E�HP�u��A�u�ЍE�P�q������   ^��]� ��U����VW�}��@(W�@p�Ѕ�t9����΋P(�GP�Bp�Ѕ�t"����΋P(�GP�Bp�Ѕ�t_�   ^]� _3�^]� ���U����VW�}��@(W�@t�Ѕ�t9����΋P(�GP�Bt�Ѕ�t"����΋P(�GP�Bt�Ѕ�t_�   ^]� _3�^]� ���U����SVW�@(��}W�@p�Ѕ���   ����΋P(�GP�Bp�Ѕ���   ����΋P(�GP�Bp�Ѕ�to����_S�΋@(�@p�Ѕ�tX����΋P(�CP�Bp�Ѕ�tA����΋P(�CP�Bp�Ѕ�t*�G��P������t�G$��P������t_^�   []� _^3�[]� �����U����SVW�@(��}W�@t�Ѕ���   ����΋P(�GP�Bt�Ѕ���   ����΋P(�GP�Bt�Ѕ�to����_S�΋@(�@t�Ѕ�tX����΋P(�CP�Bt�Ѕ�tA����΋P(�CP�Bt�Ѕ�t*�G0��P�-�����t�GH��P������t_^�   []� _^3�[]� �����U�����@(�@8]�����������������U�����@(�@<]�����������������U�����@(�@@]�����������������U�����@(�@D]�����������������U�����@(�@H]�����������������U�����@(�@L]�����������������U�����EQ�$�@(�@P��]� �U�������E�@(�$�@T��]� ���������������U�����u�u�@(�@|��]� ������U������ �@$VW�u�@���M�Q�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�Ѓ��E���P�L   ������E�P�I�I�у���_^��]� �����������U�����} �P(�����E�B8]����U��Q���VW���M�@j �@d�Ћ��h��h�  �p�IV���   �ыȃ�����M���u�@(��j��@4��_3�^��]� �@j VQ�M�@h�С����V�@(�@H�Ѕ�t�����V�u��@(�@ �Ѕ�t�   �3��E�P�t�������_^��]� �������U����VW�}��@(Q��@P�$�Ѕ�tG����GQ���$�@(�@P�Ѕ�t)����GQ���$�@(�@P�Ѕ�t_�   ^]� _3�^]� ������������U����VW�}���@(����@T�$�Ѕ�tK������G�΋@(�$�@T�Ѕ�t+������G�΋@(�$�@T�Ѕ�t_�   ^]� _3�^]� ������U����VW�}��@(Q��@P�$�Ѕ���   ����GQ���$�@(�@P�Ѕ���   ����GQ���$�@(�@P�Ѕ���   ����GQ���$�@(�@P�Ѕ�te����GQ���$�@(�@P�Ѕ�tG����GQ���$�@(�@P�Ѕ�t)�G��P�.�����t�G$��P������t_�   ^]� _3�^]� ��������U����VW�}���@(����@T�$�Ѕ���   ������G�΋@(�$�@T�Ѕ���   ������G�΋@(�$�@T�Ѕ���   ������G�΋@(�$�@T�Ѕ�ti������G �΋@(�$�@T�Ѕ�tI������G(�΋@(�$�@T�Ѕ�t)�G0��P������t�GH��P������t_�   ^]� _3�^]� �����������̡���@(� ������U����V�u�@(�6�@�Ѓ��    ^]���������������U�����@(���   ]��������������U�����@(�@]����������������̡���@(�@�����U����V�u�@(�6�@�Ѓ��    ^]���������������U�����u�u�@,Q�@�Ѓ�]� �̡���@,�@����̡���@,�@����̡���@,�@����̡���@,�@ ����̡���@,�@(����̡���@,�@$�����U�����@,�@]�����������������U�����U���@,VWR�@�Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у���_^��]� ����̡��j j �@,� �Ѓ��������������U����V�u�@,�6�@�Ѓ��    ^]��������������̡���@,�@4����̡���@,�@8�����U�����U���@,VWR�@<�Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у���_^��]� �����U�����U����@,VW�u�@@R�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]� ̡���@,�@,�����U����V�u�@,�6�@0�Ѓ��    ^]���������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����u�u�@�@\��]� ������U�����u�u�@��  ��]� ���U�������E�@�$�@ ��]� ���������������U�����EQ�$�@�@$��]� �U�������E�@�$�@(��]� ���������������U�����@�@,]�����������������U�����@�@0]�����������������U�����@�@4]�����������������U�����@�@8]�����������������U�����@�@<]�����������������U�����@�@@]�����������������U�����@�@D]�����������������U�����@�@H]�����������������U�����@�@L]�����������������U�����@�@P]�����������������U�����@���   ]��������������U�����uQ�@��  �Ѓ�]� ��U�����@�@T]�����������������U�����@�@X]�����������������U��U��u3�]� ���RQ�@ �@(�Ѓ��   ]� �����U�����@���   ]��������������U�����@�@`]�����������������U�����@�@d]�����������������U�����@�@h]�����������������U�����@�@l]�����������������U�����@�@p]�����������������U�����@�@t]�����������������U�����@���   ]��������������U�����@��  ]��������������U�����@�@x]�����������������U�����@�@|]�����������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����uQ�@��  �Ѓ�]� ��U�����@���   ]��������������U�����@���   ]��������������U��U��t���RQ�@ �@$�Ѓ���t	�   ]� 3�]� �U����Q�u�@ �u�@L�Ѓ�]� ��U�����@���   ]�������������̡���@���   ��U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]�������������̡���@���   ��U�����@���   ]�������������̡���@���   �����@���   �����@���   �����@���   �����@���   ��U����V�uV�@���   �Ѓ��    ^]�������������U�����@� ]�����@�@�����U�����@���   ]��������������U�����@��   ]��������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����@�@]�����������������U�����@���  ]��������������U�����@�@]�����������������U����E�V�u��P��������M�Q�@$�@�Ѓ���t]����M�jQ�@�@�Ѓ���u�E�P��������t3���jV�@�@�Ѓ���u���V�@�@�Ѓ���t�   �3�����H$�E�P�IH�ы���E�P�I�I�у���^��]��������U�����@�@ ]�����������������U�����@�@(]�����������������U�����@��  ]��������������U�����@��   ]��������������U�����@��  ]��������������U�����@��  ]��������������U�����M���@VWQ�@$�Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у���_^��]��������U�����M���@VWQ���  �Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у���_^��]�����U��j�u�  �E��]������������U���<����E�    SVW��t�EĻ   P��������-����M�Q�   �@�@�С���M�Q�@$�@D�Ѓ��}����uV�@�@�С��V�@$�@D�С��VW�@$�@L�Ѓ���t(����M�Q����@$�@H�С���M�Q�@�@�Ѓ���t&����H$�E�P�IH�ы���E�P�I�I�у�_��^[��]������U�����M���@VW�u���  Q�Ћ�����}W�I�I�ы��W�A$�@D�С��WV�@$�@L�С���H$�E�P�IH�ы���E�P�I�I�у� ��_^��]��U�����@��D  ]��������������U�����@��H  ]��������������U�����@��L  ]��������������U�����M����@VW�u���  �uQ�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]��������������U�����@���  ]��������������U�����@���  ]�������������̡��Vj j��@��@�Ћ�^���������U����Vj �u�@��@�Ћ�^]� �U����V�u��@j��@�Ћ�^]� ̡���@�@�����U����Vj ��M�@j V���   �Ћ�^]� �����������U�����uQ�@�@�Ѓ�]� �����U�����uQ�@�@�Ѓ����@]� U����h#  �u�@�u�@l��]� �U����hF  �u�@�u�@l��]� �U�����u�@�@t�Ћ��P���   �@X�Ѓ�]� ����U�����u�@�@t�Ћ�����uR���   �@`�Ѓ�]� ���������������U�����u�@���   �Ћȅ�u]� ���Q���   �@�Ѓ�]� ��������U�����@���   ]���������������A    ���    �A    �A   ���U�����u�u�@@�uQ�@�Ѓ�]� ���������������U�����uQ�@@�@�Ѓ�]� �����U�����u�u�@@Q�@�Ѓ�]� ��U�����uQ�@@�@ �Ѓ�]� �����U�������   �@]��������������U�������   �@]��������������U�������   �@ ]�������������̡�����   �@$��U�������   ���   ]�����������U�������   ��D  ]�����������U�����uQ�@@�@L�Ѓ�]� ����̡��Q�@@�@H�Ѓ����������������U�������   ���   ]�����������U�������   ���   ]����������̡��Q�@H���   �Ѓ�������������U��V��M��t2����U���   ��t�@@R��^]� �U�@D��tR��^]� V��^]� �����������̡���@@�@0�����U��V�u���t���Q�@@�@�Ѓ��    ^]����������U����V��V�@@�@�ЋЃ��E��t��#��С��RV�@@�@�Ѓ�^]� �U���u �E��������   �$�u�u���   �u�u��]� ����������U�������   ���   ]����������̡��Q�@H���   �Ѓ�������������U�����uQ�@H��d  �Ѓ�]� �̡���@@�@T�����U�����@@�@X]�����������������U�����@@�@\]����������������̡���@@�@`�����U�����@@�@d]�����������������U�����@@�@h]�����������������U�����@@�@l]�����������������U�����@@�@p]����������������̡���@@�@t����̡���@@�@x�����U�����@@�@|]����������������̡���@@���   ��U�����@@���   ]�������������̡���@@���   �������   �@t��U�����@@���   ]��������������U�����@@���   ]��������������U�����@@���   ]��������������U�����@@���   ]��������������U�����@@���   ]��������������U�����@@���   ]��������������U�����@@���   ]��������������U��V�u���t���Q�@@�@�Ѓ��    ^]���������̡���@@�@0�����U�����MjQj �@@�@4�Ѓ�]����U�����MjQh   @�@@�@4�Ѓ�]�U�����u�u�@@j �@4�Ѓ�]���̡���@|� ������U��V�u���t���Q�@|�@�Ѓ��    ^]���������̡���@|�@ �����U��V�u���t���Q�@|�@(�Ѓ��    ^]����������U�����@ �@H]�����������������U��}qF uGW�}��t>������u���   �@D�С���u�@@�@,�Ћ�����ЋA��W�u�@p��_]������������U�����@��T  ]��������������U����SVW�@@�u�@,�Ћ�����u�I@�I,�ы�������y��h��hE  ����Ph��hE  ������P��T  �Ѓ�_^[]�����̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������3�� �����������3�� �����������U��M�E�A4�E�A �E��E�A0�E�A ��A8c��A<h��A@���AD���AHr��ALm��AP|��Al���AX���A\��A`���Ad���ATw��Ah���Ap��At���A(�A,    ]��������������U���   h�   ��`���j P�� j �u��`����u�u�uP�����E h�   �E���`���P�u�uj��  ��8��]�����U���   V����	  �����   S�u�M����������M�Q�@�@�С���M�j j�hp��@Q�@�Ѓ��E��M�P����j j��E�P�E�P��d���P������P�E�P�������P�E�P��������P�  ���M���������M��������d���������M����������M�Q�@�@�Ѓ��M�������[t	V�	  ����^��]� ������U��V�u���r  �����^]� ������Q��  YË�`��`$��`(��`,��`4��`8��`@��`3���������������U��E�     3�]� �������������̋�PP�   ����U����   V�u��u3�^��]�h�   ��@���j P�� �E����@����΍�@�����`���ǅD��� �h�   P��u�E�h��E����E����E�m��E�r��PPj��  ��^��]�U��j�u���������u]Ë�]�b����̡���@��   ��U����V�u�@�6��$  �Ѓ��    ^]������������U����V��V�@�u��(  �Ѓ���^]� ������������U����Q�u�@��,  �Ѓ�]� ��U����Q�u�@��,  �Ѓ����@]� �������������U��E��t�P�3ҡ��RQ�@��8  �Ѓ�]� ������U�����uQ�@��<  �Ѓ�]� ��U�����u�u�@�uQ��@  �Ѓ�]� ������������U�����u�u�@Q��D  �Ѓ�]� ���������������U�����uQ�@��H  �Ѓ�]� ��U�������@VW�u��L  Q�M�Q�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]� ������������̡��Q�@��T  �Ѓ������������̡��Q�@��P  �Ѓ�������������U�����uQ�@��X  �Ѓ�]� ��U�����uQ�@��l  �Ѓ�]� �̡���@��0  �����@��4  �����@��p  �����@��t  �����@��\  ��U����V�u�@�6��`  �Ѓ��    ^]������������U���u����u�u�@�u�u��d  Q�Ѓ�]� ������U���u����u�u�@�u�u��h  Q�Ѓ�]� �����̡��Q�@�@�Ѓ����������������U���u����u�u�@�uQ�@X�Ѓ�]� ������������U�����uQ�@�@\�Ѓ�]� ����̡��Q�@�@ ��Y�U�������@Vh�  Q���   �M�Q�Ћ��P���   �@8�Ћ�����E�P���   �	�у���^��]��������������U�����@��   ]��������������U�����u�u�@�uQ�@�Ѓ�]� ���������������U���u����u�u�@�uQ���   �Ѓ�]� ���������U�����@�@$]�����������������U���u����u�u�@�uQ�@(�Ѓ�]� ������������U���u����u�u�@�uQ�@,�Ѓ�]� ������������U���u(����u$�u �@�u�u�@`�u�u�u�uQ�Ѓ�(]�$ �������������U����VW���@W�@�Ћ����W�J�I���u���H�u�u�Q�N�QPj �B4j W�Ѓ�(_^]� ���������������U���u ����u�u�@�u�u�@4�u�uQ�Ѓ� ]� ���U�����u�u�@Q�@@�Ѓ�]� ��U�����uQ�@�@D�Ѓ�]� ����̡��Q�@�@L�Ѓ���������������̡��Q�@�@L�Ѓ���������������̡��Q�@�@P�Ѓ����������������U�����uQ�@�@T�Ѓ�]� �����U�����uQ�@�@T�Ѓ�]� ����̡��Q�@�@h�Ѓ����������������U�����u�u�@Q���   �Ѓ�]� ���������������U�������@V�u�u���   Q�M�Q�Ћuj PV�    �F    ������   �I�ы���E�P���   �	�у� ��^��]� ��������̡���@� ������U����V�u�@�6�@�Ѓ��    ^]���������������U���u����u�u�@�u�u���   Q�Ѓ�]� ������U����V�u�@�6�@�Ѓ��    ^]���������������U��QVW�}�����n ���V�@�@h�Ѓ������u"�@h��h�  ��0  �Ѓ�_3�^��]� �M��E    �@Q�MQ�u���   V�Ѓ���tыM�3���~�d$ �E����tP����l �M�F;�|�EP�}������   _^��]� �������������U��QVW�}����n ���V�@�@h�Ѓ������u"�@h��h�  ��0  �Ѓ�_3�^��]� �M��E    �@Q�MQ�u���   V�Ѓ���tу} t�3�9u�~2�E����t"���Q�@�@h�Ѓ���t�E���4���k F;u�|΍EP襼�����   _^��]� �����U�����@��x  ]�������������̡���@��|  ����Q�@���   �Ѓ�������������U�����uQ�@���   �Ѓ�]� �̡���@���   ��U����V�u�@�6���   �Ѓ��    ^]������������VW���O�����W����G �G0�G@�GP�    �G`    �Gd    �Gh    �Gp�Gx�����G|   _^�����������V���X   �N^�O������������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7��������xP t$V������j j j�pP�ˍGP�ݿ���H ���^�    �` t����w`�@�@�Ѓ��G`    _[�������������h��h�   h�h�   �7�������t������3��������U��V�uW�>��t���K����O�C���W�ݷ����_�    ^]�U����SVW�@��W��   �_dS�wx�w`�uV�Ѓ��G|����   �? ��   �; ��   �wpV�_hS�u��  ����u&�W�����h��h  �@��0  �Ѓ��u�O�P������觾���xP u����"��蕾��j j j�pP�ˍGP聾���H ��ЉG|��t���[����G|_^[]� �G|�Gx����_^[]� �G|�����    ����6�@�@�Ѓ��    �G|_^[]� �V������W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������U��QW���d �G`t~S�];_xttV�7�ΉE�u�跽���xP u����#��襽���M�S�u�pPj�GP落���H ��ЉG|^��u�E�_x��t�    �G`[_��]� �M�Gx������t�3�[_��]� �����������U��E��t	�Ap� �yd t�Ah]� 3��y|��]� ���U���u ����u�u�@�u�u�@�u�uQ�Ѓ� ]� ���U�����uQ�@�@�Ѓ�]� ����̡��Q�@�@��Y�U�����u�u�@Q�@�Ѓ�]� �̡���@� ������U����V�u�@�6�@�Ѓ��    ^]���������������U��VW���D����u���u�x@�u�1����H ���_^]� ����U��VW�������u���u�xD�u�����H ���_^]� ����W�������xH u3�_�V���ֻ���ύpH�̻���H �^_�����U��W��赻���xL u3�_]� V��蠻���u���u�pL�u荻���H ���^_]� U��W���u����xP u���_]� V���_����u���u�pP�u�u�I����H ���^_]� ������������U��W���%����xT u���_]� V�������u���u�pT������H ���^_]� ��U��W�������xX u���_]� V���Ϻ���u�ύpX�º���H ���^_]� �����U���SVW�}�م�t.�M�������菺���ˍpL�E�P聺���H ��ЍM��@����u��tW����M�Q�@�@�С���M�VQ�@�@�С���M�Q�@�@�Ѓ����+����H@��t���VQ�@�@�Ѓ�_^[��]� ���������U��VW��������u�΍xH�����H ���_^]� ����������U��W���Ź���x` u
� }  _]� V��譹���u�ύp`蠹���H ���^_]� ���U��SVW��胹���x` u� }  �#���o����ύp`�E���P�\����H ��Ћ�����]S�I�I�у�;�>���S�@�@�Ѓ�;�)�������u���u�pDS�u�
����H ���_^[]� _^�����[]� U��W�������xP u
�����_]� V���͸���u���u�pP�u�u�u�u豸���H ���^_]� ����U��W��蕸���xT u
�����_]� V���}����u���u�pT�m����H ���^_]� U��W���U����xX tV���G����u�ύpX�:����H ���^_]� �������������U����E��E�    P�u�E�    �E�    �E�    �E�    �E�    �f ����t(�M��t!�u�����u��u��@�u�Q�@X�Ѓ���]�3���]��������������������������������U��M�]�`����U��M�]�`����V��h �Vh���$��F    ���h���@P� �Ѓ��F��^����������̃y �$�u����q�@P�@��Y���U��I��u3�]� ���j �u�@P�uQ�@�Ѓ�]� ���U��I��t����uQ�@P�@�Ѓ�]� ��������������U��I��t����uQ�@P�@�Ѓ�]� ���������������    ���A    �V����t&���Q�@P�@L�С���6�@P�@<�Ѓ��    ^����������������U��SVW�����t���Q�@P�@<�Ѓ��    �G    �M�]h ��O���Sh��h���@PQ�u�@8��3����9u~E���x u�@   ����HP���p�A�Ѓ����V�7�@P�@@�Ћ���F�A;u|�3�9_^��[]� �����������U���u�E�u�p�,���]� ��������U��SVW��3�9w~=�]���V�7�@P�@@�ЋЃ���t-���j Sj�APR�@�Ѓ���tF;w|�_^�   []� ����7�@P�@L�Ѓ�3�_^[]� ������������̡���1�@P�@D�Ѓ��������������̡���1�@P�@H��Y���������������̡���1�@P�@L��Y���������������̡���@P�@P�����U�����@P�@T]����������������̡���@P���   ��U�����@P���   ]��������������U��M�]�`����U��V��~ �$�u����v�@P�@�Ѓ��Et	V�_�������^]� ������8����A    �A    �A    ���V��~ �8�u����v�@4� �Ѓ��F    �F    ^���������������̸   ����������̸   �����������3�� ������������ �������������U����V��h�  �@4�v�@$���u����u�u�@4�u�v�@�Ѓ�2�^]� ���������������U���u��u�u�u�P]� ��������3�� ����������̸   � ��������� �������������U��Q���SVW�@�ً}3��ω]��@ ��=INIb�  ��   =SACbmt)=$'  t
=MicM�f  ���W�P$�   _��^[��]� ��MQ�M��u�Q�ˉu�P��t����u�u��@4�s�@�Ѓ��   _��^[��]� =ARDb�  �����j j�@���   �Ћ؋ϡ��j j�@���   �ЋM�����j j�@���   �ЋM����j j�@���   ���u�M�PVW�S�R�   _��^[��]� ����P�   _��^[��]� =NIVb_tF=NPIbt.=ISIbuV�3���  P���r  P���V�   _��^[��]� ���W�P_^[��]� ����P�   _��^[��]� =cnyst_��^[��]� �����j hIicM�@���   �Ћ��WP�R _^[��]� �������U���,V��~ t~����v�@4�@�Ѓ} t���P�F�I0�p�Al�Ѓ�^��]� ���E��M��E�    hARDb������NP�E�P�E�P�q  ����M�Q���   � �Ѓ��M������^��]� ������������U�����u�q�@4�@l�Ѓ��   ]� �������������̡���q�@4�@�Ѓ�������������̡���q�@4�@�Ѓ�������������̡���q�@4�@�Ѓ�������������̡���q�@4�@|�Ѓ�������������̡���q�@4���   �Ѓ�����������U�����u�q�@4�@(�Ѓ�]� ���U���u����u�u�@4�q�@,�Ѓ�]� �������������U�����u�u�@4�q�@0�Ѓ�]� ����q�@4�@4��Y���������������U�����u�q�@4���   �Ѓ�]� U�����u�q�@4�@ �Ѓ�]� ���U�����u�q�@4�@$�Ѓ�]� ���U����V�uW���   ��V�@�Ѓ������V���   u �@@�Ћ��P�w�I4�A �Ѓ�_^]� �@�Ѓ������u'���   V�@8�Ћ��P�w�I4�A$�Ѓ�_^]� �@h4�h  ��0  �Ѓ�_^]� ����������U�����u�u�@4�q�@D�Ѓ�]� U�����u�u�@4�q�@H�Ѓ�]� U�����u�u�@4�q�@L�Ѓ�]� U�����u�u�@4�q�@P�Ѓ�]� U����SVW���   �ً}W�@�Ѓ���������   �@��   �uV�Ѓ������V���   u6�@@�Ћ����W���   �I@�ы��VP�s�I4�AP�Ѓ�_^[]� �@�Ѓ������u=���   V�@8�Ћ����W���   �I@�ы��VP�s�I4�AH�Ѓ�_^[]� h4�h�  ��   W�Ѓ��������   ���   �uV�@�Ѓ������V���   u6�@@�Ћ����W���   �I8�ы��VP�s�I4�AL�Ѓ�_^[]� �@�Ѓ������u=���   V�@8�Ћ����W���   �I8�ы��VP�s�I4�AD�Ѓ�_^[]� h4�h�  �
h4�h�  �@��0  �Ѓ�_^[]� �����U���u����u�u�@0�u�q���   �Ѓ�]� �������U���u����u�u�@4�u�q�@�Ѓ�]� ����������U���u����u�u�@4�u�q�@�Ѓ�]� ����������U���u,����u(�u$�@4�u �u�@T�u�u�u�u�u�q�Ѓ�,]�( ��������U���u����u�u�@4�u�q��  �Ѓ�]� �������U����h����h����h�����u�@4�uh�����@Th����h����h�����u�q�Ѓ�,]� ����������U�����u�q�@4�@8�Ѓ�]� ���U�����u�q�@4�@<�Ѓ�]� ���U�����u�u�@4�q���   �Ѓ�]� ������������̡���q�@4�@@�Ѓ�������������̡���q�@4��  �Ѓ�����������U�������E�@4�$�q��  �Ѓ�]� ������U���u����u�u�@4�u�q�@X�Ѓ�]� ���������̡���q�@4�@`��Y��������������̡���q�@4�@d�Ѓ��������������U���u����u�u�@4�u�q��   �Ѓ�]� �������U���u����u�u�@4�u�u�@\�u�q�Ѓ�]� ����U�����u�u�@4�q��  �Ѓ�]� �������������U�����u�u�@4�q�@h�Ѓ�]� U�����u�u�@4�q��  �Ѓ�]� �������������U�����u�u�@4�q�@p�Ѓ�]� U���V��M�hYALf�
������P�v�R4�Bl�Ѓ��M��-���^��]���������U��QVW�}�M���t����Mj j�@���   �Љ�u��t����Mj j�@���   �Љ����M�VW�@4�q�@p�Ѓ�_^��]� �������U���u����u�I�u�@0�q���   �Ѓ�]� �������U���u����u�u�@4�u�q�@x�Ѓ�]� ����������U�����u�q�@4�@t�Ѓ�]� ���U���u����u�u�@4�u�u���   �q�Ѓ�]� ����U���u����u�u�@4�u�u���   �q�Ѓ�]� ����U������S�E�    �ًM�E�    �@W�{j ���   j�ЋM�E����j j�@���   �ЉE��M����Q�M�Q�@0�w�@`�С���s�@4�@�Ћ���U�j R�U�I0R�U�R�U�RP�C�p�Ah�Ѓ�,�} _[t(�} t(�M�U�;�~<�E��;�}3�M��U�;�~)�E���} u�M�U�;�~�E��;�}�   ��]� 3���]� ���U���u�E������@4�D$�E�$�u���   �q�Ѓ�]� �����U���u����u�u�@4�q���   �Ѓ�]� ���������̡���q�@4���   �Ѓ�����������V��Vh�M�h�����@0� �Ѓ��F�F    ��^�����V��N�h���t���Q�@0�@�Ѓ��F    ^������̸   ����������̸   ����������̸   � ��������3�� �����������3���������������� �����������������������������U����VW�}��@�ϋ@ ��=NIVb��   ��   =TCAbwtM=$'  t3=MicM��   �����j hIicM�@���   �Ћ��WP�R_^]� ���W�P_�   ^]� �����j hdiem�@���   �Ћ��WP�R_^]� =INIbu�~ u�����F   �P_^]� �~ t�����P_^]� =atni@t1=ckhct=ytsdu;����P_�F    3�^]� ����P_^]� 襭  _3�^]� =cnys����_3�^]� ����������U��V��N��u3�^]� ���j j j �@0j j �u ���   j �ujQ���u����u�u�@0�uj �u���   �v�Ѓ�D^]� ����������̋I��u3�á��Q�@0�@�Ѓ�����̋I��u3�� ���Q�@0�@�Ѓ�� U���V�q��u�E�p�    ^��]� �E�H����Q�u�M��@0RVQ���   �Ћuj PV�    �F    ������   �I�ы���E�P���   �	�у�$��^��]� ��������U�����u�q�@0���   �Ѓ�]� ����q�@0���   �Ѓ����������̡��j j j �@0j j j ���   j j j4�q�Ѓ�(�������̡��j j j �@0j j j ���   j j j;�q�Ѓ�(��������U�����u�q�@0�@�Ѓ�]� ���U��I��t'���j j j �@0j j j �u���   j jQ�Ѓ�(]� �����������U���u����u�u�@4�q�@,�Ѓ�]� �������������U�����u�u�@4�q�@0�Ѓ�]� ����q�@4�@4��Y���������������U��V�q��u3�^]� �E�H����Q�u�@0RV�@�Ѓ�^]� �����������U��V�q��u3�^]� �E�H����QRV�@0���   �Ѓ�^]� �����������U��E3�h���h  �P��j ��BRj �u�u�   ]� ���U���$VW���M�htniv�y�������M��uhulav�@�@4�С���M�hgnlfhtmrf�@�@4�С���M��uhinim�@�@4�С���M��uhixam�@�@4�С���M��uhpets�@�@4�С���M��uhsirt�@�@4�ЋM �u$��  �u�����t,���Qh2nim�M܋@�@4�С���M�Vh2xam�@�@4�ЍE܋�P�u�E�P�S������P���   �@8�Ћ�����E�P���   �	�у��M�����_��^��]�  ������U���$V��M�htlfv�:�������M��E���@�$hulav�@,�С���M��u,htmrf�@�@4�С���M��E���@�$hinim�@,�С���M��E���@�$hixam�@,�С���M��E$���@�$hpets�@,�С���M��uDhsirt�@�@4���U0W�f.џ��Dz�E8f.����D{?����M܃��@�$h2nim�@,�С���M��E8���@�$h2xam�@,�С���M��u@hdauq�@�@4�ЍE܋�P�u�E�P�������P���   �@8�Ћ�����E�P���   �	�у��M�������^��]�@ ������������U���u,W�j ��$htemf�E$�� �D$�E�D$�E�D$�E�$�u����]�( ���������������U���Mf.�����%h����D{�Y��^��Uf.�����D{�Y��^��u,W�j ��$hrgdf�E$�� �Y��^��D$�E�L$�T$�$�u�o���]�( �����������U���u,�X�W�j ��$htcpf�E$�� �^��D$�E�^��D$�E�^��D$�E�$�u�����]�( �����������U���0�E�M���u����@���   �Ѕ�u��]� SVW���,�  htlfv�MЋ�������u�����fn���ɋy��Y��E��E��$�n� �]��F�$�`� �E�M��]��^E�G,�$hulav�С���M�hmrffhtmrf�@�@4�Ћu�����fn���ɋx��Y��E��E��$��� �]��F�$�� �E�M��]��^E�G,�$hinim�Ћu�����fn���ɋx��Y��E��E��$螘 �]��F�$萘 �]��E�M��^E�G,�$hixam�С���M�������@�$hpets�@,�С���M�j hdauq�@�@4�С���M�Shspff�@�@4�С���M��u hsirt�@�@4�ЋM��E�P�u�E�P�������P���   �@8�Ћ�����E�P���   �	�у��M��a���_��^[��]� ������U���$V��M�hCITb���������M��uhCITb�@�@8�С���M��uhsirt�@�@4�С���M��uhulav�@�@4�ЍE܋�P�u�E�P�`������P���   �@8�Ћ�����E�P���   �	�у��M�譾����^��]� ����U��V�q��u3�^]� �E�E�H����Q�u �@0���@(�D$�E�$�uRV�Ѓ�$^]� U����E�Vj �u��MP����P�u�������������E�P�I�I�у���^��]� �����������U��V�q��u3�^]� �E�H����Q�MQ�@0RV�@,�ЋM3҃�9U�^]� �������������U��V�q��u3�^]� �E�H����Q�u�@0RV�@,�Ѓ�^]� �����������U��V�q��u3�^]� �E�H����Q�u�@0RV�@0�Ѓ�^]� �����������U��VW���O����   �E�P�0���R�u�@0VQ�@0�Ѓ���tf� t`�E�H����Q�p0�E��P�F0R�w�Ѓ���t8���t1�E�H����Q�p0�E��P�F0RW�Ѓ���t_�   ^]� _3�^]� ��������������U��QV�q��u	3�^��]� �EW�E�    �H����Q�M�Q�@0RV�@8�Ћ�����t:�U���t3����uR�A�@�Ћu�����t���V�@�@��V�Ǎ������_^��]� ����������U��V�q��u3�^]� �E�H����Q�u�@0�uR�@<V�Ѓ�^]� ��������U��E��V���u����@���   �Ѕ�u^��]� W���]�  �v����t!�E�H����Q�M�Q�@0RV�@0�Ѓ���fnǍM�������Y���D$�E��Y���$�E _�o �E� ��^��]� �����������U�������@V��M�Q�@�Ѓ��E���P�u�U�������t�M�E�P�ӗ������E�P�I�I�у���^��]� �����U��V�q��u3�^]� �E�H����Qj j �@0j j j ���   j Rj1V�Ѓ�(^]� �������������U����Vj �u�@��M���   ��h���h  �j j jj P�u���E���^]� U����Vj �u�@��M���   ���u$���u j �u�u�uP�u����^]�  �U������W�V����M�@�$�u���   ���E8��j �u@�]����D$�E0�$�u,�E$�� �D$�E�D$�E�D$�E��$�u����^��]�< ����U������W�V����M�@�$�u���   ��j j ��W��]���$htemf�E$�� �D$�E�D$�E�D$�E��$�u�8���^��]�$ �U������W�V����M�@�$�u���   ���Uf.�����%h���]���D{�Y��^��Mf.�����D{�Y��^�j j ��W���$hrgdf�E$�� �Y��^��D$�E��T$�L$�$�u�t���^��]�$ �������������U������W�V����M�@�$�u���   ���X�W�j j �����]�$htcpf�E$�� �^��D$�E�^��D$�E�^��D$�E��$�u�����^��]�$ �������������U���0���(��V��M�Q�ufE��@�M�Q�M���   ��j �u ���u�o �E��u�E�P�u�u�x���^��]� �U������0�@VW���M��@Q�С���M����@Q�u�MЋ��   Q�M�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�Ѓ��E����uj P�u����������E�P�I�I�ы���A�M�Q�@�Ѓ���_^��]� ���U���dV��M��O�������MP�u�R�E�P���   ��P�M��ڑ���M�����j j �E�P�M�蒒��P�u������������E�P�I�I�у��M��ؑ���M��Б����^��]� �������U���P����U�E�V�uW�����t+�����W��΋@�$R���   ���]��E��E�����M�W�Q�ufE��M��E��@Q�΋��   �Ћw�o �E��~@f�E؅�u
_3�^��]� �E�E�H����Q�u �Mȋ@0���@(�D$�E��$QRV�Ѓ�$_^��]� ���U��V�q3���t)�E�H����Q�MQ�@0RV�@,�Ћ���3�9E�����P�u�Q�M�R0�ҋ�^]� ��������������U��V�q��t!�E�H����Q�MQ�@0RV�@,�Ѓ�������u�u�A�M�@4�Ћ�^]� ������U���V�q��t!�E�H����Q�M�Q�@0RV�@0�Ѓ���������E��A�M�$�u�@,�Ћ�^��]� �������U���(���E�VP�ufE��u�����������E�P�u�Q�M�R@�ҋ�^��]� �����������U���V��W�WfE�~�E�����   �E�H����Q�M�Q�@0RW�@0�Ѓ���tx�~��tq�E�H����Q�M�Q�@0RW�@0�Ѓ���tN�v��tG�E�H����Q�M�Q�@0RV�@0�Ѓ���t$����M�Q�u�M�@�@H��_�   ^��]� _3�^��]� ���������U�������@V��M�Q�@�Ѓ��E���P�u�����������E�P�u�Q�M�R8�ҡ���M�Q�@�@�Ѓ���^��]� ��������������U���,V��M��?�������M�Q�@�@�Ѓ��E���P�u�m�������u����M�Q�@�@�Ѓ�� �E�P�M��Վ������M�Q�@�@�Ѓ�����M�P�E�P�u�R<�ҍM�貍����^��]� ���������U��� V�qW��E�fE���t%�E�H����Q�M�Q�@0�M�QRV�@<�Ѓ����U���t����A�M�Q�MR�@H�ЋU���t������E��M�@�$R�@,�Ћ�^��]� ���U��E3�Vh���h  ��8�p�   ��RE�3���j ��@Pj V�u�����^]� ��������������U���u �U3��u�:��P�u�u�u�r�u����]� ���U��U3��E4�:��P�u<���D$�E,�$�u(�E �� �D$�E�D$�E�D$�B�$�u�}���]�8 ���������U��E3�W��8�H��Rj ��$htemf�E �� �D$�E�D$�E�D$�$�u����]�  ������U��E3��U���%h��8�h��f.�����D{�Y��^��Mf.�����D{�Y��^�Rj ��W�$hrgdf�E �� �Y��^��D$�T$�L$�,$�u�v���]�  ��U��E3��X�W��8�P��Rj ��$htcpf�E �� �^��D$�E�^��D$�E�^��D$�$�u����]�  ��U��U3��:��P�u�B�u�uP�u�u�����]� �����U��E3��u�8��RP�u�����]� ��������������U���$V��M�hgnrs�ڭ���E�M��E�����E�   Qj�@�M܋��   �С���M�Q���   � �ЋE�M��E�������E�   Q�@�M�j���   �С���M�Q���   � �Ѓ��E܋�P�u�E�P�������P���   �@8�Ћ�����E�P���   �	�у��M��]�����^��]� ����U��W�y��u3�_]� �E�EV�H����Q�u �p0���E���D$�E�$P�F(RW�Ѓ�$^_]� ���������̡��j j j �@0j j j ���   j j j �q�Ѓ�(��������U��I��u3�]� ����u�u�@4Q��  �Ѓ�]� ��U��I��u3�]� ����u�u�@4Q�@h�Ѓ�]� �����U��I��u3�]� ����u�u�@4Q�@p�Ѓ�]� �����U��I��u3�]� ����u�u�@4Q��  �Ѓ�]� ��U���u����u�u�@0�u�q���   �Ѓ�]� �������U�����P0�E�pj j j �u�uj �0���   j=�q�Ѓ�(]� �����������U�����P0�E�p�uj j j��uj �0���   j=�q�Ѓ�(]� �����������U��E�x��u��EС���2�@0�u�q�@@�Ѓ�]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u�u���   �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u�u���   �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   �u�ujQ�ЋE���(��]� ���������������U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �uj*Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�uj �u���   j	Q�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�uj �u���   j
Q�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u�u���   �uj'Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u�u���   �uj,Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �uj:Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j j �u�E�    �u�@0j j j)���   Q�ЋE���(��]� ���U��Q�I��u3���]� ����U�Rj j �u�E�    �@0j �u���   j j j)Q�ЋE���(��]� ���U��I��u3�]� ���j j j �u�@0�u�u���   j �ujQ�Ѓ�(]� ��U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u�u���   j �uj>Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U����j j j �u�@0�u�u���   j �uj.�q�Ѓ�(]� �������������U��V�q��u3�^]� �E�H����Qj j �@0j j �u���   �uRjV�Ѓ�(^]� �����������U��V�q��u3�^]� �E�H����Qj j �@0j j j ���   j RjV�Ѓ�(^]� �������������U��V�q��u3�^]� �E�H����Q�u�@0RV�@\�Ѓ�^]� �����������U���SVW�u�ٍM���{���EP�E�P�M��
|����tj�}�I �M��tI���Q���   �@H�ЋS������tN�w���j j j �A0j �u����   V�7jR�Ѓ�(��t"�EP�E�P�M��{����u�_^�   [��]� _^3�[��]� ���U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U����VW�}��@4�w� �ЋE�G    �w�H����Q�u�@0WR�v���   �Ѓ��G3Ʌ���_��^]� �������U��I��u3�]� ���j j j �u�@0�u�u���   j �uj/Q�Ѓ�(]� ��U��U��u3�]� �r�B    ����u�q�@0���   �Ѓ�]� ���������U��I��u3�]� ���j j j �@0j j �u���   j j jQ�Ѓ�(]� ����̡��j j j �@0j j j ���   j j j6�q�Ѓ�(��������U��I��u3�]� ����u�u�@0�uQ�@D�Ѓ�]� ��U��I��u3�]� �u����u�u�@0�u�u�@H�uQ�Ѓ�]� ��������̋I��u3�á��Q�@0�@X�Ѓ������U��I��u3�]� ����u�u�@0Q�@L�Ѓ�]� �����U��Q��u3�]� ����H0�E   �P�APR�Ѓ�]� ��U��I��u3�]� ����uQ�@0�@P�Ѓ�]� ��������U��I��u3�]� �u����u�u�@0�uQ�@T�Ѓ�]� ���������������U���VW���M��N����E�M�P�0���RQj �@0j j j ���   j Vj8�w�Ћ���(��t�M�E�P�|����M��d���_��^��]� ����������U��EV�P�0���R�u�@0j j j ���   j j Vj9�q�Ѓ�(^]� ��������U��EV�P�0���R�u�u�@0�u�u�@hV�q�Ѓ�^]� ��������������U��QVW�}�M���t����Mj j�@���   �Љ�u��t����Mj j�@���   �Љ����M�VW�@0�q�@`�Ѓ�_^��]� �������U���u����u�u�@0�q���   �Ѓ�]� ����������U�����U�@0��t*���   R�q�Ћ�����uR�A0���   �Ѓ�]� �u�@|�q�Ѓ�]� ��U���u����u�u�@0�u�u�@p�q�Ѓ�]� �������U���u����u�u�@0�u�u�@d�q�Ѓ�]� �������U����j j �u�@0�u�u���   �uj �uj3�q�Ѓ�(]� ������������U��Ej j j ����j j j �@0j Rj�q���   �Ѓ�(]� �������������U��Ej j j ����j j j�@0j Rj�q���   �Ѓ�(]� �������������U��Ej j j ����j j j �@0j Rj�q���   �Ѓ�(]� �������������U��EV�P�0���Rj j �@0j j j ���   j Vj"�q�Ѓ�(^]� ���������U��EV�P�0���Rj j �@0j j j ���   j Vj5�q�Ѓ�(^]� ���������U��EV�P�0���Rj j �@0j j �u���   j Vj<�q�Ѓ�(^]� ��������U����Vj j �@0��j j j �u���   j �uj�v�С���u�v�@0�@t�Ѓ�0^]� �������̡��j j j �@0j j j ���   j j j�q�Ѓ�(��������U����j j j �@0j j j �u���   j j�q�Ѓ�(]� ���j j j �@0j j j ���   j j j�q�Ѓ�(��������U����j j j �@0j j j ���   j �uj�q�Ѓ�(]� U����j j j �@0j j j �u���   �uj&�q�Ѓ�(]� ��������������̡��j j j �@0j j j ���   j j j(�q�Ѓ�(�������̡��j j j �@0j j j ���   j j j#�q�Ѓ�(��������U����j j j �@0j �u�u���   j �uj+�q�Ѓ�(]� �������������̡��j j j �@0j j j ���   j j j0�q�Ѓ�(��������U�����u�q�@0���   �Ѓ�]� U���V�u ��M��L�������M��uh8kds�@�@4�С���M Q�M��E     Q�@0j �u�u���   �u�u�uj2�v�Ћu �M��(������^��]� �������̡���q�@0���   �Ѓ�����������U��I��u3�]� ���j j j �@0j j j ���   j �uj-Q�Ѓ�(]� �����U������Wj ���M�@j���   �ЋM�E����j j�@���   �ЉE��M����Q�M�Q�@0�w�@`�С���U��H0�E�pR�U�R�U�R�U�R�0�Ah�w�Ѓ�(�} _t(�} t(�M��U�;�~<�E��;�}3�M��U�;�~)�E���} u�M��U�;�~�E��;�}�   ��]� 3���]� �����U��SV�uW��u�q����]��j hdiuM�@���   �Ћ���tI;>u	_^3�[]� �����j hIicM�@���   ��;�u�����j h1icM�@���   �Шu��>_^�   []� ���������U������(�@V�u��hfnic�@T�ЋЅ�t���j
�A�ʋ��   �Ѕ���   ����M�hfnicQ�΋@�@P��P�M�讖���M��Ɩ���u�E�P���Ȗ���M�谖������΋@�@ �Ѓ��t����΋@�@ �Ѕ�u�����hfnic�@�@$�С�����uj
�@�@8��^��]������������̡���q�@0���   �Ѓ�����������U���$V��M�hmnrs�ڕ������M��uj�@�@4�ЍE܋�P�u�E�P�s������P���   �@8�Ћ�����E�P���   �	�у��M��������^��]� �������U���$�DSSS�} V��SSSSE��M�P�M�������M܋@�@ �Ћ��jP�Q�M܋B4�ЍE܋�P�u�E�P��������P���   �@8�Ћ�����E�P���   �	�у��M��$�����^��]� �����������V��Vh�M�h�����@0� �Ѓ��F�F    ������F   �F    ^�V��N�h���t���Q�@0�@�Ѓ��F    ^�������U��V��N�F    ��tg���j j j �@0j j j ���   j j jQ���u����u�u�H03�9E�u����
j P�v���   �Ѓ�D��t�~ t
�   ^]� 3�^]� ��������������U��E�A�I��u3�]� ���Q�@0�@�Ѓ�]� �����U����S�]V�@��ˋ@ ��=ckhc��   t|=cksatb=TCAb��   �����Wj hdiem�@���   �Ћ��SW���F   �R�~ ��t��t��u3��΃���P�J���_^��[]� �~ ti����P^[]� �~ tV���j j j �@0j j j ���   j j j �v�Ѓ�(��t*�F    �   ^[]� =atnit�u��S�x���^[]� ^3�[]� ����������U��Q�y �M���   S�]V�uW�}��wp�$�(;9u��   �^9u��   �S9u��   �H9u��   �=�E;�~6;���   �,�E;�|%;�~}��E;�|;�|p��E;�~;�~c�9uu\���j j j �@0j j j ���   j �uj�q�Ѓ�(fn����j���D$fn�����$S��x  �E����@    _^[��]� �Y:d:o:z:�:�:�:�:�:����U��W��� �6  V�u����   �$��<�Ef/E�  �   �Ef/E��   �   �Mf/M��   �   �Mf/M��   �|�Uf/Uvp�E f/���   �_�Uf/UrS�E f/���   �B�Uf/Ur6�E f/�w�)�Uf/Uv�E f/�sf��Ef.E���DzT���j j j �@0j j j ���   j �uj�w���E ��(�u(���D$�E�$V�uw  ���G    ^_]�$ �t;�;�;�;�;�;�;<1<U���E j���D$�E�D$�E�$�u�u�]���]�  ���������U���E j���D$�E�D$�E�$�u�u����]�  ���������U���E j���D$�E�D$�E�$�u�u�����]�  ���������V��Vh�M�h�����@0� �Ѓ��F�F    ������F   ^��������V��N�h���t���Q�@0�@�Ѓ��F    ^�������U����V��M�@�@ ��=cksat]=ckhct�u���u�o���^]� j j j j j �F   ���j j j �@0j �v���   �Ѓ�(��t#�F    �   ^]� �~ t����P^]� 3�^]� �������������U��V��Vh�M�h�����@0� �ЋM���F�E�F    �F   ����F���j hmyal�@���   �ЉF��t��t�F    ����Mj
hhfed�@���   �ЉF��^]� U����V��M�@�@ ��=ytsdt�u���u����^]� ����v�@0���   �Ћ�����P�   ^]� ����������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U���V�u�V�E�    �    �B    ���������E�    j ���   �E�PR�I�ы���E�P���   �	�у���^��]� ����������̋A��uË ���������������������U��V���PD��t�E9Ft
�F�΋�PH^]� ���������̋A�������������U��j0�u�l  ��]���������������U��j0�u�C�  ��P�l  ��]������U����E�j0�u�uP�I�  ��P�`l  ����M�Q�@�@�Ѓ���]���������U����E�j0�u�u�uP�f�  ��P�l  ����M�Q�@�@�Ѓ���]������U��j$�u��k  3Ƀ�������]�����U��j$�u胼  ��P��k  3Ƀ�������]������������U����E�Sj$�u�uP�x�  ��P�k  ���3ۃ��E�P�ËI�I�у���[��]������������U����E�Sj$�u�u�uP腽  ��P�<k  ���3ۃ��E�P�ËI�I�у���[��]���������U�����u�u�@j ���   �Ѓ�]�U�����u�u�@�uj ���   �Ѓ�]��������������U�����@���  ]��������������U�����@0���   ]��������������U�����M����@0VW�u���   �uQ�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]��������������U���4���SV�u�@WV�@�С�����M3ۋ@SS���   �ЋM�E����Sj�@���   �Ћ����M  3ɉM�d$ ��~k����M�Q�@�@�С���M�j j�ht��@Q�@�С�����΋@�@<�ЋȍU���j�j�R�@Q�΋@L�С���M�Q�@�@�Ѓ�����M�W�u��@0Q���   �Ћ��Mܡ��Q�@�@�С���M�QW�@�@�С���M�Q�@�@�С�����΋@�@<�ЋȍUܡ��j�j�R�@Q�΋@L�С���M�Q�@�@�С�����MC��
�M�@j Q�M���   �ЋM�E�A���j Q�M�P���   �ҋ��������_��^[��]����U�����@0���   ]��������������U�����@0���   ]��������������U�����@0���   ]�������������̋�W�R�J��A(�P$j j h����?l  �������������̸x������������U���(V��M�WQ�΋�P(�V����t&���j j j �A0j j j ���   Wj jR�Ѓ�(����M�Q�@�@�С���M�Q�@�@�ЋN����t����U�j Rj �@0jj?j �@HQ�Ѓ�����M�Q�@�@�С���M�Q�@�@�ЋN����u3��:����U�Rj j j h  
 j�U��E�    �@0Rh�  j���   Q�Ћ}���(����M�Q�@�@�Ѓ���u_3�^��]á���M�Q�@�@�ЋN����t����U�j Rj �@0j j8j �@HQ�Ѓ�����M�Q�@�@�ЋN����t���jQ�@0�@P�Ѓ�����M�Q�@�@�Ѓ��M��C���Ph   h  K j;�E��Ph	��h�  ��������M�Q�@�@�Ѓ��M��e����N��t���Q�@0�@X�Ѓ��N��t���Q�@0�@X�Ѓ��N��t&���j j j �@0j j j���   j j jQ�Ѓ�(j�v$��d  ���   _^��]�U���V��Wj�N�,����F4    W��F8    �F<    �F(���h�   �v�@0�@�С���M�Q�@�@�С���M�j j�h���@Q�@�Ѓ��E��  �E��E�    ��j j P�E�P��������M�Q�@�@�Ѓ��Nj j�[���_^��]������U���\���VW���Mȋ@Q�@�С���M�j j�h���@Q�@���G(�YX�����E��  �E�    �@�,ȋ@(Q�M�Q�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M��8�@�@<�Ћ��j�j��Q�M�QP�M�BL��j j �E��P�E�P���������M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ��M�htats詂������M�jj�@�@0�С���M��G(���@�$j�@,�ЍE��E��  P�E��E�    P�E���P��������M�Q���   � �Ѓ��4 t_����O0�@P�@h�ЋG4��t�w8�Ѓ��G<�G8    �G4    ����h4�h�  �@��0  �Ѓ�����O0�@P�@l�ЍM�����_^��]� ����������U������@�@V�uW�@ ������=MicMtG=fnic��   j�M�舁���MP�ρ���M�跁������Mjj�@�@4��_�   ^��]� �����j hIicM�@���   ��=���uhtats�M��)�������M�j j�@�@0�ЍE��E��  P�E��E�    P�E��P贸������M�Q���   � �Ѓ��M������O�G   ��t���Q�@0�@�Ѓ��u��V����_^��]� ����U��mV��t3�^]� j�N����j�`  �N���F    ��t���Q�@0�@�Ѓ��   ^]� j���֢��j�`  ��3�����������U���E�A(]� ��������������̍A�������������U��VW��~4 t@�I ���h4�hs  �@��0  ��j
��k  ����v �@P�@�Ѓ���uM9F4uá���N0�@P�@h�Ѓ~4 t:���h4�h�  �@��0  �С���N0���@P�@l���r���_3�^]� �E�N0�F8�E�F4���S�@P�@l�Ѓ~4 t#j
�ik  ����v �@P�@�Ѓ���u99F4uݡ���N0�@P�@h�Ћ~<�N0�F<    ����RP�Rl��[��_^]� [_3�^]� U����M�V�~���M�����t �@4Q�@�Ѓ���t$��M�Q�u���R(�1�@0�u�@�Ћȃ���u�M�3���~����^��]Ë�U�R�u�P ���M����@�@ �Ѓ��t����H0�E�P�u�Ix�у��M��~~����^��]��������U����Vj �u�@��M���   �Ћ���u�    �F^]� ��u9Ft�   ^]� ���������U��V�uW��;uuz����Mj htsem�@���   �Ѕ�u\����Mj hrdem�@���   �Ѕ�u>�E�E�H��t1����Uj RV�@0Q�@,�Ѓ���t�u���  _�   ^]� _3�^]� ���������������U������@�@VW���M��@Q�С���M�Q�@�@�С���MЃ��@Q�u�M����   Q�M�Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�С������@V�@�С���M�VQ�@�@�Ѓ����%  ����M�Q�@�@�Ѓ�_^��]� ���������U���SV�u��;u��   ����Mj htsem�@���   �Ѕ���   ����Mj hrdem�@���   �Ѕ���   ����M�Q�@�@�ЋM�E���u��E�    P�E�P�h�����u3��4�������@V�@�С���M�VQ�@�@�Ѓ����A  �   ����E�P�I�I�у���^[��]� ^3�[��]� ���U����Vj �u�@��M���   �Ћ���u�    �F^]� ��u9Ft�   ^]� ���������U���V�uW��;uup����Mj htsem�@���   �Ѕ�uR����Mj hrdem�@���   �Ѕ�u4�M�E�E��EP�E��u�P�ɼ����t�u���  _�   ^��]� _3�^��]� ����U������W�V����M�@�$�u���   �Ћ�]����u�E��    �F^��]� ��u�Ff.E����D{�   ^��]� ����U���SV�u��;u��   ����Mj htsem�@���   �Ѕ�um����Mj hrdem�@���   �Ѕ�uO�EW��E��H��t=����U�j RV�@0Q�@0�Ѓ���t!�E������$�,  ^�   [��]� ^3�[��]� �����U���H���W�V���E��M�Q�ufE�@�M�Q�M���   ���o �~H��EЃ��u�F�    f�N^��]� ��u5�Ff.EП��Dz�Ff.E؟��Dz�Ff.����D{�   ^��]� U���4�ES�]�M�V�uW�};�t;�t;���   ����Mj htsem�@���   �Ѕ���   ����Mj hrdem�@���   �Ѕ�ui�MW��E��E��E�E�P�E��E�P�E�u�P�E�}�PfẺ]�������t.�oE̋M������ �~E�f�@��  �   _^[��]� _^3�[��]� ����U��� ���(��V��M�Q�ufE��@�M�Q�M���   ���o ��E����u�    �F^��]� ��u�E�P�FP��   ����t�   ^��]� ������U���SV�u��;u��   ����Mj htsem�@���   �Ѕ�ui����Mj hrdem�@���   �Ѕ�uK(���M�E��E�P�u�E��u�PfE��Y�����t"�oE���ˋ�� �0  �   ^[��]� ^3�[��]� ���������U���V�uW�}�f.���Dz�Ff.G���D{Y�G���Y��E��E��$��N �F�Y�]��E��E��$��N �E����]�f.E����D{_�   ^��]�_3�^��]����U��V��N�h���t���Q�@0�@�Ѓ��E�F    t	V��G������^]� ���������������U��V��~ �8�u����v�@4� �Ѓ��E�F    �F    t	V�rG������^]� ��������U�����u�E�    �A]� ��u�A;Et�   ]� U�����u�E�    �A]� ��u�Af.E���D{�   ]� ����U�����u�oE�    �A�~Ef�A]� ��u6�Af.E���Dz �Af.E���Dz�Af.E���D{�   ]� ����������U��V�����u�oE�    �F^]� ��u�EP�FP��������t�   ^]� �����������U��V�����u �    ����P�FP�EP�B�Ѓ��"��u����MQ�N�@�@x�Ѕ�t�   ����MQ�@�@�Ѓ�^]� ��������U�����@ �@h]�����������������U����V�u�@@�6�@�Ѓ��    ^]���������������U�����uQ�@ �@�Ѓ�]� �����U�����uQ�@ �@�Ѓ�]� ����̡��Q�@ �@��Y�U��VW�}�����r�����WV�J �I�у���_^]� ����U�����uQ�@ �@ �Ѓ�]� ����̡��Q�@ �@,�Ѓ���������������̡��Q�@ �@0�Ѓ����������������U�����uQ�@ �@4�Ѓ�]� ����̡���@ � ������U��V�u���t���Q�@ �@�Ѓ��    ^]����������U������� V��W�}��~D�F<    �F8    �F@    �FH    �FL   �FP    �FT    ����   �E��P��5  P�N��Q���M��"N������8  �F�ύE�P�-A  W�o �F����@@�@,�Ћ�����tH���j h6  �Q�ϋ��   �҉FP�ϡ��j h5  �@���   ��_�FT^��]� �F   _^��]� ������������̋I@��t���Q�@�@D�Ѓ�ø   �̡���@���   ��U����V�u�@�6���   �Ѓ��    ^]�����������̡��Q�@���   ��Y��������������U��EWɋMW�HH H0H@HP� (���@(��f�H�@0f�H(W�f�H@����@Hf�HX�o� �~Af�@]�������U��EWɋMW�HH H0H@HP� (���@(���@0f�H(W�f�H@f�H����@Hf�HX��@�A�@8�A�@X]������������U���W�W�V�uNN N0N@NP�(���F(���F0W�f�Nf�N(f�N@����FH�Ef�NX��3 �E��E��C �U�f(�fWP����VX�N@�FP�V8^��]�����U���W�W�V�uNN N0N@NP�(���F(���F0W�f�Nf�N(f�N@����FH�Ef�NX�/3 �E��E� C �U�f(�fWP����V�NH�F(�VX^��]�����U���W�W�V�uNN N0N@NP�(���F(���F0W�f�Nf�N(f�N@����FH�Ef�NX�2 �E��E�pB �M����F0fWP��N�F �N8^��]���������U������   V�u�V �F(��^(�Y��Y��X�(��Y��X���C f(�W�f.џ��Dz2W�fD$X(��D$P�D$h�D$`�D$8�D$X�D$�K����^��N�Y��L$�L$X�N �Y��L$8�L$`�N(�Y��L$P�L$h�N0�^8(��V@�Y�(��Y��X�(��Y��X��C f(�W�f.џ��Dz#W��L$0f�$�   ��$�   �D$@�E����^��N0�Y��L$@��$�   �N8�Y���$�   �N@�Y��L$0�fP�VH(��^X(��Y��Y��X�(��Y��X��iB f(�W�f.џ��Dz$W��L$fD$x��$�   f(��L$x�<����^��NH�^P�VX�Y��Y��Y��L$x��$�   �T$�E��$�   �\$p�L$H����  �$��h�D$0��fWP��$�'  ���\$�D$��/ fWP�fT@�f/��v6�D$h݄$�   ��O �\$ ݄$�   ݄$�   ��O �\$(�D$(��  �D$`W��D$X�D$�O �D$0f/���\$ ��  �(��\D$ �D$ �  �D$@���$�I&  ���\$(�D$(�D$�/ fT@�f/��vR�D$0fWP��D$�D$݄$�   �%O �T$HfWP��\$�T$�D$�D$X� O �\$ �  �D$hW��D$�D$8fWP��D$�D$��N W�f/D$@�\$ ��  ���\D$ �D$ �  ��(�fWP��$�_%  ���\$ �D$ �-. fT@�f/��v6݄$�   �D$X�UN �\$(݄$�   ݄$�   �>N �D$(�\$�C  W��D$�D$8fWP��D$�D$݄$�   �N W�f/D$H�\$�	  �D$fWP��D$��  �D$8��fWP��$�$  ���\$(�D$(�D$�Y- fWP�fT@�f/��v-�D$h�D$X�|M �\$ ݄$�   ݄$�   �eM �\$�v  �D$xW�݄$�   �D$ �CM �D$8f/���\$�E  �D$�X��D$�,  �D$P���$��#  ���\$ �D$ �, fT@�f/��vB�D$8fWP��D$�D$�D$X�L �D$0fWP��\$(�D$�D$�O����T$HW�fWP�݄$�   �T$�D$�D$�lL W�f/D$P�\$�s  �D$�\��D$�Z  ���$�	#  ���\$�D$��+ fT@�f/��vE�T$HfWP��T$�D$݄$�   ��K �D$8fWP��\$ �D$�D$�����݄$�   W��D$X�D$�K W�f/D$p�\$ ��  �D$ fWP��D$ �  (��Y�f(��Y��X���< ���f(�f/��l$@��   �T$8W��\$P�Y�f(��Y��L$�XT$�X�f/��r�L$�5���f/�r���D$�(��t" �\$PW��D$�d$pf/�v���f/�����f/��D$ ��  �(��\D$�D$�  �\$W�f/����T$H�L$�^�v^f/��r���fWP��   ���f/�r���fWP��l(��<J �l$@f(�fWP�W��Mf/��r
����5���f/�r
����(���I ��f(��l$@W��X�f/��T$�T$0v�X(��T$0�T$�d$p�^�(��0& �D$ �D$0�/) �D$@�D$0�9 �\$@W��L$8�Y\$�YD$P�Y��X��X�f/��rf(��#���f/�r
���(��  W��D$�L$8f/�v�(��\�f(��D$�E�oD$^�L$� f�H��]ÍI pa4bcze�c�d����U������V�uW�W�}��W�F(��Y�(��Y��X���9 ���f(�f/��T$v<�GW�f/���v(���f�N_^��]�(���f�N_^��]��Gf/����^�vTf/��r���fWP��z���f/�r���fWP��Z(���G �T$fWP��Bf/��r
����&���f/�r
����(��G �T$�X���G�^��$ �F��W�_�F^��]�������������U���   V�uW��f.��E���D��   �Ff.����Dzq�Ff.����Dzb�EW�^HH H0H@HP� (���@(���@0f�HW�f�H(f�H@����@Hf�HX��]��E�W�}�;6 ��u7�E���(& �E��F�6 f(��F�M��& �E��5f(���M���% �E��F��5 �E��F��% �E��F��5 �E��F�% f(���p������  �$� q�m�E��e�f(��YU�f(�P�}�f(��YǍE�Pf(��YߍE��Y��Y��\�f(��Y��M�f(��X��Y��Y��U��U�f(��YE��E�f(��Ye��Y��\��E�f(��Y��Y��]��E�f(��YE��U��X��M��  �m�f(��YE�f(��YU�f(��}�fWP��E�f(��YE�f(��YM��Ye��Y��X��m��E��YE��M�(��YM��\��U��E�f(��Y��E�f(��Y�fWP��E�f(��Y��YU��Y��X��   �e�f(��E�f(��m��M��}��Y��Y�fWP��E�f(��Y��E�f(��Y��E�f(��Y�f(��Y��Y��E�f(��Y��X�f(��Y��M�f(��\��Y�f(��Y��Y��U��Y��X��Yu��E�P�\��eЍE�P�u��E��M��  �e؍E��m�f(��}�f(��Y�f(�P�YE��E�P�YߍE�f(�fW%P��YM��YU��e��\�f(��Y��M�f(��YM��E�f(��YE��X�f(��Ym��U��U��Y��Y��X�f(��Y��\��M��E�f(��YE��Y��]��E��u���   �}��E��e�f(��YU�f(�P�m�E��Y�f(�P�Y]��E�f(��Y��Y��\�f(��Y��M�f(��X��Y�(��Y��U��U��Y��Y��E�(��Y��Y��X�f(��Y�fW%P��Y��\��M��e��u��E��E��E�fW-P��m��MW�P��x����]�W�Pf�x����4  �E_^��]��e�f(��YM�(ċE�YE�f(�_�m���p���f(��YM�f(�^fWP��Yu��Y]��E��YU�f(��YE��Ym��Y}��X���p���(��\�f(��Ye��YM�f(��YE��Y]�f��\��E��YE��X�W�fWP�XX X0X@XP�E�W�� �E�f��oE��H�M�f��p0�@Hf�Xf�P(f�h@f�xX��]Ë��k�lMm�on�n��������U�������   V�uW�o�o^ �oV��$�   �oF0f���$�   �oF@f(���$�   �oFP�Y���$�   f(��Y��T$ (�f��X�f(�)T$P�Y��X��1 W�f.����Dz)W��L$PfD$ �D$(�D$�D$ �D$8�7����^�f(��YD$ �D$8f(��YF �YL$P�D$�L$P��$�   ��$�   (��Y���$�   �Y��X�(��Y��X���0 W�f.����Dz,W�fD$ (��D$�D$(�D$@�D$ �D$ �A����^�f(��Y�$�   �D$ f(��Y�$�   �Y�$�   �D$@�L$��$�   ��$�   (��Y���$�   �Y��X�(��Y��X��80 f(�W�f.ʟ��Dz)W�f(�fD$h�D$p�d$h�D$H����9���f(��^�f(�f(��Y�$�   �Y�$�   �Y�$�   �l$H�L$@�XL$8�d$�X��\��Y��f/�s$���f/�r
���(��} f(��L$�\L$H�\$�\\$P�u�}f(��L$�Y���T$�\T$ �(��Y��\$�^�T$�X��V(��Y��X��/ W�f.����Dz	W�f(��<����^��D$�d$�Y��Y��D$h�D$�d$p�Y�fT$h�f�F�f.����Dz2�Ff.����Dz#�Ff.����Dz(���f�N�_^��]��������U���������@W�W�V�uW�}NN N0N@NP�(���F(���F0W�f�N�FHf�N(f�N@f�VX�f.����Dz"�Gf.����Dz�Gf.����D��  �Ef.����D��  �Y���E��+ �D$�E� ��_�D$�G�Y��Y��\$�X�f(��Y��X��V- f(�W�f.˟��DzW�fD$0�|$8�t$0�'����^��7��\$�Y��Y��Y��D$�l$�Y��Y��Y����f(��Y�f(��Y��\$�Y�f(��Y��|$f(��Y��D$(f(��Y�f(��Y��D$(��Y�f(��Y�(��Y�(�����D$ �D$�Y��Y|$�L$0�XL$�D$�X��Xt$ �\�(��\��X�f�����Vf�N(�L$�XL$ �\�(��\L$(�X|$(f��oD$0�n0�\D$f�N@����\�f��FHf�NX_��^��]���������U���p�EV�uW�o�E���wB�$�${����F�X��X��\V�=���Ff(��\�X�����f(��\F�X��V�XӋ}���]�f��M��\�U��^(��]��E��$�]��&- �M؃��(��]��\M��Y�f/�f(��M��X�U�r�\��\��M��U��M����\O�^��M��E��$�M��, �M����(��]��\M��Y�f/�f(��M��XW�U�r�\��\��M��U��W���~N�\��^��M��E��$�M��A, �MЃ��(��]��\M��Y�f/�f(��M��XW�U�r�\��\��M��U��]����\�^��]��E��$�]���+ �M���(��]��\M��Y�f/�f(��M��X�U�r�\��\��M��U��U����\W�^��U��E��$�U��a+ �E����(��]��\E��Y�f/�f(��E��XW�U�r�\��\��E��U��E����\G�^��E��E��$�E���* �M����(��]��\M��Y�f/�f(��Xg_^r�\��\��@��]�fT��U�fT؋EfT��X��]�fT��X��M�fT��X��]�fT��X�f/�v�oE�� f�`��]��oE�� �E�f�@��]��w�w�w�w�w�w����U����M�Q�	(��Y�Y��Y��X�(��Y��X�W�f.��M����Dz�E �@��]ËU�E�B�p�8�\���j�\��`f(��\̋E�Y���Y��Y�X�(��Y��I�X���^U��Y��Y��Y��X���X��X��\��\�� �B�\��h�@��]�������������U��E�M�p�f(��yf(��!�X�i�Y̋E�Y��X�f(��Y��X��Y���Y��Y��Y��\��\��\�� �x�h]����������A    ���d   �U��E�A    �]� �������������U����@i�� %����fn�������X����^���E��E���]���U����@i�� %����fn�������X����^���Y���\���E��E���]���U������V��~ �  �-��W��5���%���@i�� ���������fn�����X����Ai�� �^�%����fn�������Y��X����\��^��T$�Y��\�f(��D$�Y�(��Y��X�f/��L$�p���f.˟��D�b���f(���8 �Y���^D$��$ f(��F   �YD$�YL$�Y���N�X���D$�D$^��]��F����F    ^�����]����������������U������V��~ �  �-��W��5���%���@i�� ���������fn�����X����Ai�� �^�%����fn�������Y��X����\��^��T$�Y��\�f(��D$�Y�(��Y��X�f/��L$�p���f.˟��D�b���f(��x7 �Y���^D$�# f(��F   �YD$�YL$�Y(��N�D$�D$^��]��F�(��F    ^��]��������������U��E��Hf(�f/��pvf(�f/�vf(�f/�f(�vf(�f/�vf(�W�f/���   f(��=���^��\����f/�v�E�h ]�f.�f(��\ş��Dz
�\��^��2f.˟��Dz(��\��^��X����\��^��X�(��^ �f/�v�X���E��x�X]ËE�` ]�������������U�������V�uf/F��Vv(�(���   f.�����DzW��Y ����M��E��$�M���# �m����~�%���]��M�f(��\��V�,�f(�f(��Y��\�H�Y��\�f(��\��Y��Y��\��Y��w>�$�D�f(�f(��4f(�f(�(��+f(�f(��!(�f(��(�f(�f(��(�f(�f(ӋE^��@�P��]ÍI �� �
���������̡���@���   ��U����V�u�@�6���   �Ѓ��    ^]������������U����j �u�@���  �Ѓ�]����U����V�u�@�6���  �Ѓ��    ^]������������U�����@���   ]��������������U����V�u�@�6���   �Ѓ��    ^]������������U��� ���W�j j j fE��E�    �E��E�    �H�E�Pj �E�P�EPPP�u��d  �u�u�uj �Ѓ�8��]�����U�����uQ�@���   �Ѓ�]� ��U���u����u�u�@�u�u���   �uQ�Ѓ�]� ���U���u����u�u�@�u�u���   �uQ�Ѓ�]� ���U���u����u�u�@�uQ���   �Ѓ�]� ���������U���u����u�u�@�uQ��  �Ѓ�]� ���������U�����u�u�@Q���   �Ѓ�]� ���������������U��VW�}�����G�����WV�J���   �у���_^]� �U�����uQ�@���   �Ѓ�]� ��U�����uQ�@��  �Ѓ�]� �̡��Q�@��0  �Ѓ�������������U�����u�u�@Q��t  �Ѓ�]� ���������������U���u����u�u�@�uQ���  �Ѓ�]� ���������U��U��tA���    t8�MV��  ;q}(��t	�E�    �	��  �t	�E�    ^]�����    ����������V����t���Q�@��<  �Ѓ��    ^������������U��V����t���Q�@��<  �Ѓ��    ����u�u�@�u��8  ��3ɉ��������^]� ��������������V����t���Q�@��<  �Ѓ��    ^������������U��	��t����u�u�@Q���  �Ѓ�]� ���������U��	��t����u�u�@Q���  �Ѓ�]� ���������U�����@��P  ]��������������U�����@��T  ]��������������U�����@��X  ]��������������U���V�u����\E�^(��E��E��$�E�� �M����(��]��\M��Y�f/�f(��M��XE�r�\��\��M���E�^��]�������������U��EW�AA A0A@AP�o ��~@�Ef�A�o �A�~@�Ef�A(�o �A0�~@�Ef�A@�o �AH�~@��f�AX]� ������U���Mf/��r���]����f/�r���]�(��) �E�E]��������������̡��Q�@L���   �Ѓ�������������U�����u�u�@LQ���   �Ѓ�]� ���������������U����V��V�@L���   �Ћȃ������u�@LQ�u���   V�Ѓ�^]� ���   �@P�Ћ��P���   �M�BH��^]� �������������̡��Q�@L��(  �Ѓ�������������U�����u�u�@LQ��,  �Ѓ�]� ��������������̡���@L� ������U����V�u�@@�6�@�Ѓ��    ^]��������������̡���@L���   ��U����V�u�@@�6�@�Ѓ��    ^]���������������U�������u�@LQ�M�Q�@�ЋM��P�IB���M��aB���E��]� ��������U�����u�u�@LQ�@�Ѓ�]� ��U�����uQ�@L���   �Ѓ�]� �̡��Q�@L�@�Ѓ���������������̡��Q�@L�@�Ѓ���������������̡��Q�@L�@�Ѓ����������������U�����u�u�@L�uQ�@ �Ѓ�]� ���������������U�����uQ�@L��4  �Ѓ�]� ��U�����u�u�@L�uQ�@$�Ѓ�]� ���������������U���u����u�u�@L�uQ�@(�Ѓ�]� �����������̡��Q�@L�@,�Ѓ���������������̡��Q�@L�@0�Ѓ���������������̡��Q�@L�@4�Ѓ���������������̡��j Q�@L�@8�Ѓ��������������U�����u�u�@LQ��  �Ѓ�]� ���������������U�����@L���   ]��������������U�����@L���   ]��������������U�����@L��l  ]��������������U�����@L���   ]��������������U�����@L���   ]��������������U�����@L���   ]��������������U�����@L���   ]��������������U�����@L���   ]��������������U�����@L���   ]��������������U�����uQ�@L�@<�Ѓ�]� �����U�����@L���   ]�������������̡��Q�@L�@��Y�U�����u�u�@LQ�@@�Ѓ�]� ��U����j �u�@LQ�@D�Ѓ�]� ���U����j�u�@LQ�@D�Ѓ�]� ���U����j �u�@LQ�@H�Ѓ�]� ���U����j�u�@LQ�@H�Ѓ�]� ��̡��Q�@L���   �Ѓ�������������U�������u�@LQ�M�Q��  �ЋM��P��=���M���=���E��]� �����U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ���  j �E܋�P�E�P��?�����M����i�  ��t3������M�Q���   �@8�Ѓ�������E�P���   �	�у���^[��]����������U���$V�E��E�   ���E�   P�M��E��  �E�    �E�    �X�  j�E܋�P�E�P�w?���M��φ  ����M�Q���   � �Ѓ�^��]�����U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ��  j �E܋�P�E�P��>�����M����Y�  ��t
�M���� ����M�Q���   �@L�ЋM��P�+������E�P���   �	�ыE��^[��]� ���������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �7�  j �E܋�P�E�P�6>�����M���詅  ��t
�M����� ����M�Q���   �@L�ЋM��P�{������E�P���   �	�ыE��^[��]� ���������U���$����E�    �E�    V���   ���u�M�Q�@(�Ѓ��E��  �E��E�    �M��E�    P�n�  j�E܋�P�E�P�=���M���  ����M�Q���   � �Ѓ�^��]� ��������U���$����E�    �E�    V���   ���u�M�Q�@(�Ѓ��E��  �E��E�    �M��E�    P�ނ  j�E܋�P�E�P��<���M��U�  ����M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �g�  j �E܋�P�E�P�f<�����M����ك  ^��[tW��E��E������M�Q���   �@<�Ѓ�����M�Q�]����   � ���E�����]����������������U����E�E�V���E�   P�M�E��E��  �E�    �E�    赁  j�E��P�EP��;���M�,�  ����M�Q���   � �Ѓ�^��]� ���������������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �7�  j �E܋�P�E�P�6;�����M���詂  ��t3������M�Q���   �@8�Ѓ�������E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    虀  j�E܋�P�E�P�:���M���  ����M�Q���   � �Ѓ�^��]� ���U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �'�  j �E܋�P�E�P�&:�����M���虁  ��t8����E܋uW�P���   �����F�	�у���^[��]� ����M�Q���   �@P�Ћ���u�o ���   �E�P��	�у���^[��]� �������������U���$����E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�.  j�E܋�P�E�P�M9���M�襀  ����M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �~  j �E܋�P�E�P�8�����M����)�  ��t8����E܋uW�P���   �����F�	�у���^[��]� ����M�Q���   �@P�Ћ���u�o ���   �E�P��	�у���^[��]� �������������U���$����E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�}  j�E܋�P�E�P��7���M��5  ����M�Q���   � �Ѓ�^��]� ��������U�������@Lj�u���   Q�M�Q�Ѓ��o �E� ��]� ������������U�������@Lj �u���   Q�M�Q�Ѓ��o �E� ��]� ������������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ��|  j �E܋�P�E�P��6�����M����9~  ��t8����E܋uW�P���   �����F�	�у���^[��]� ����M�Q���   �@P�Ћ���u�o ���   �E�P��	�у���^[��]� �������������U���$����E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P��{  j�E܋�P�E�P��5���M��E}  ����M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �W{  j �E܋�P�E�P�V5�����M�����|  ��t8����E܋uW�P���   �����F�	�у���^[��]� ����M�Q���   �@P�Ћ���u�o ���   �E�P��	�у���^[��]� �������������U���$����E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�^z  j�E܋�P�E�P�}4���M���{  ����M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ��y  j �E܋�P�E�P��3�����M����Y{  ��t3������M�Q���   �@8�Ѓ�������E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    �Iy  j�E܋�P�E�P�h3���M���z  ����M�Q���   � �Ѓ�^��]� ���U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ��x  j �E܋�P�E�P��2�����M����Iz  ��t8����E܋uW�P���   �����F�	�у���^[��]� ����M�Q���   �@P�Ћ���u�o ���   �E�P��	�у���^[��]� �������������U���$����E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P��w  j�E܋�P�E�P��1���M��Uy  ����M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �gw  j �E܋�P�E�P�f1�����M�����x  ��t3������M�Q���   �@8�Ѓ�������E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    ��v  j�E܋�P�E�P��0���M��@x  ����M�Q���   � �Ѓ�^��]� ���U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �Wv  j �E܋�P�E�P�V0�����M�����w  ��t3������M�Q���   �@8�Ѓ�������E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    �u  j�E܋�P�E�P��/���M��0w  ����M�Q���   � �Ѓ�^��]� ����������t��t��t3�ø   ���̡��Q�@L�@L�Ѓ���������������̡��Q�@L�@P�Ѓ����������������U�����u�u�@LQ�@T�Ѓ�]� ��U�����uQ�@L��  �Ѓ�]� ��U�����uQ�@L���   �Ѓ�]� �̡��Q�@L�@X�Ѓ����������������U�����u�u�@L�uQ�@\�Ѓ�]� ���������������U������0�@LSV��@�Ћ؅�u^[��]� W�M��+���u�E��E�    �E؍M����E�    �E�    �E�    �E�    �]Ћ@h]  �@0�С����j j S���   �@�Ѕ���   ���S�@L�@�Ћ�������   �d$ ������   �΋R(�ҋ��uԍE�Ph�   �  ����tq�M��tj���j ���   ���   �ЋЅ�tO���V���   �ʋ@<�С���M�Q���   ���   �Ѓ���t���V�@@�@�Ѓ������d����*���S�@@�@�С���M�Q���   ���   �Ѓ�3ۍM��p  �M��*��_^��[��]� ������������̡��Q�@L�@`�Ѓ���������������̡��Q�@L�@d�Ѓ����������������U�����uQ�@L�@h�Ѓ�]� ����̡��Q�@L��D  �Ѓ������������̡��Q�@L�@l�Ѓ����������������U�����uQ�@L���   �Ѓ�]� �̡���@L�@�����U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@L���   ��Y�������������̡��Q�@L���   �Ѓ�������������U���u����u�u�@L�u�u���   Q�Ѓ�]� ������U�����u�u�@L�uQ���   �Ѓ�]� ������������U���u����u�u�@L�uQ��   �Ѓ�]� ���������U�����u�u�@L�uQ��   �Ѓ�]� ������������U�����@L��H  ]�������������̡���@L��L  ��U�����@L��P  ]��������������U�����@L��T  ]��������������U�����@L��p  ]��������������U�����@L��t  ]��������������U�����@L���  ]��������������U�����@L���  ]��������������U�����@L���  ]�������������̡���@L���  ��U��U$V�u�Eh��h��h��hp�R�u �q�u�Q�u������@L�$�u���   VQ�Ѓ�4^]�  �������̡���@���   �����@���   ��U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U����V�u�@�6���   �Ѓ��    ^]������������U����V�@L�@�Ћ���u^]á��j �u�u�@�uV��h  �Ѓ���u���V�@@�@�Ѓ�3���^]������������U����j �u�H�E�� P�u��h  �u�Ѓ�]�������U�����@���   ]��������������U�����@L���   ]��������������U���u ����u�u�@�u�u���   �u�u�Ѓ�]����U��� ���W��E��E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4���jP�QL�΋��   �ЋE��E�E�Ph=���u��>
  ������   ����M�Q���   ���   �Ѓ��E�    �M��y  ��^��]���U��� ���W��E��E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4���jP�QL�΋��   �ЋE��E�E�Ph<���u��	  ������   ����M�Q���   ���   �Ѓ��E�    �M���   ��^��]���U�����@L���   ]��������������U�����@L���   ]�������������̡���@L��  �����@L��@  ��U��M�]� �����U��M�u��P]�U��M�u�u��P]��������������U���u�M�u�u��u�P]�������̡�����   �AP���   ��Y��������U�����uQ�@8�@D�Ѓ�]� ����̡���@8�@<�����U����V�u�@8�6�@@�Ѓ��    ^]���������������U���u����u�u�@8�u�u�@�uQ�Ѓ�]� ������U���u����u�u�@8�u�u�@Q�Ѓ�]� ��������̡���@8� ������U����V�u�@8�6�@�Ѓ��    ^]���������������U�����u�u�@8�uQ�@�Ѓ�]� ���������������U�����u�u�@8Q�@�Ѓ�]� �̡��Q�@8�@�Ѓ����������������U�����uQ�@8�@ �Ѓ�]� �����U���u����u�u�@8�u�u�@$Q�Ѓ�]� ���������U�����u�u�@8Q�@(�Ѓ�]� ��U�����u�u�@8�uQ�@,�Ѓ�]� ���������������U�����u�u�@8�uQ�@�Ѓ�]� ���������������U�����u�u�@8Q�@0�Ѓ�]� ��U�����u�u�@8�uQ�@4�Ѓ�]� ���������������U�����uQ�@8�@8�Ѓ�]� �����U��M����P�APP�A@P�A0P�A P�AP���   Q�u�Ѓ�]�������������̡���@���   �����@���  ��U�����@�@,]�����������������U�����@���  ]��������������U����V�uV�H�I�ы��V�I�I8�у���^]����̡���@�@<�����U�����@�@@]����������������̡���@�@D����̡���@�@H�����U�����@�@L]�����������������U�����@�@P]�����������������U�����@��<  ]��������������U�����@��,  ]��������������U���u����u�u�@�u�u���   h�2  �Ѓ�]�����U�����@�@]�����������������U�����M��� �@Q�@�С���M�j j�hD��@Q�@�С���M�Q�@�@�С���M�Q�M�Q�@�@�С���M��� �@�@<�Ћ��j�j��u�Q�M�P�BL�С���M�Q�@�@�С���M�Q�@�@�С���M�Q�@�@�Ѓ���]����U�����@���  ]��������������U�����@��8  ]��������������U�����M����@VWQ��  �Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]����U�����M����@VWQ��  �Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]����U�����@��x  ]��������������U�����@��|  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@�@T]�����������������U�����@�@X]�����������������U�����@�@\]����������������̡���@�@`�����U�����@���  ]�������������̡���@�@d����̡���@�@h�����U�����@�@l]�����������������U�����@�@p]�����������������U�����@�@t]�����������������U�����@��D  ]��������������U�����@��  ]��������������U�����@�@x]�����������������U�����@��@  ]��������������U��V�u���������V�u�I�I|�у���^]���������U�����@���   ]��������������U�����@��d  ]��������������U�����@��h  ]��������������U�����@���  ]�������������̡���@���   ��U��V�u���R�����V�I���   �у���^]��������̡���@��`  ��U�����@��  ]��������������U�����M���@�uQ���   �ЋM���o ��~@��f�A��]������U�����@���  ]��������������U���u����E���@�D$�E�$�u���   �Ѓ�]�����������U�����@���   ]��������������U�����@���   ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@��   ]��������������U�����@��  ]��������������U�����@��l  ]�������������̡���@���  ��U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����M����@VW�u���  Q�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]�U�����M����@VW�u���  Q�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]�U�����@���  ]��������������U�����@���  ]��������������U�������U�R�U�R�@�U�RQ���   �Ѓ����#E���]����������������U�������U�R�U�R�@�U�RQ���   �Ѓ����#E���]����������������U�������U�R�U�R�@�U�RQ���   �Ѓ����#E���]����������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@���   ]��������������U�����@��  ]��������������U�����@��\  ]��������������U�������u�H�E��uP��t  �у���������M��^����E��]��������U�����@��H  ]��������������U�����@��T  ]�������������̡���@��p  ��U�����@��8  ]��������������U���  ��3ŉE��EP�u������h   P��O ����x	=�  |#����h �hH  �@��0  �Ѓ��E� ���������QhH��@��4  �ЋM���3���  ��]������������������������U���u(�E�u$�u �P�u����u�u�@0�u�u���   RQ�Ѓ�(]�$ ������U���u(�E�u$�u �P�u����u�u�@0�u�u���   RQ�Ѓ�(]�$ ������U���u(����u$�u �@0�u�u���   �u�u�u�uQ�Ѓ�(]�$ ���������̡��Q�@0���   �Ѓ�������������U�����u�u�@0Q���   �Ѓ�]� ���������������U���u����u�u�@0�uQ���   �Ѓ�]� ��������̡��Q�@0���   �Ѓ�������������U���u����u�u�@0�uQ���   �Ѓ�]� ��������̡���@0���   ��U����V�u�@0�6���   �Ѓ��    ^]������������U�����M����@V�u�u��X  �uQ�Ћuj PV�    �F    ������   �I�ы���E�P���   �	�у� ��^��]����������U���4VhLGOg�M�������j P�E��IhicMCP��X  �Ћ�����E�    �E�    j ���   �M�RQ�@�С���M�Q���   � �Ѓ� �M��i������M�Q���   �@T�Ѓ���u
�M����� ����M�Q���   �@T�ЋM��P�������E�P���   �	�ыE��^��]������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����M����@VWj �u��t  �u�u�uQ�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у�(��_^��]������U�����M����@V�u�u���  �u�uQ�Ћuj PV�    �F    ������   �I�ы���E�P���   �	�у�$��^��]�������U������4�@��p  �Ѕ���   h���M��U������M��uh���@�@4�С���M��uh���@�@4�С���M�j Q�M��@hicMCQ��X  �Ћ�����E�    �E�    j ���   �M�RQ�@�С���M�Q���   � �С���M�Q���   � �Ѓ�$�M�������]����������U������4�@V��p  �Ѕ�u����uV�H�I�у���^��]�Wh!���M��\������M��uh!���@�@4�С���M�j Q�M��@hicMCQ��X  �Ћ�����E�    �E�    j ���   �M�RQ�@�С���M�Q���   � �С���M�Q���   �@H�Ћ�����}W�I�I�ы��WV�A�@�Ћ���E�P���   �	�у�4�M�������_^��]������������U������4�@V��p  �Ѕ�u����uV�H�I�у���^��]�Wh����M��<������M��uh����@�@4�С���M�j Q�M��@hicMCQ��X  �Ћ�����E�    �E�    j ���   �M�RQ�@�С���M�Q���   � �С���M�Q���   �@H�Ћ�����}W�I�I�ы��WV�A�@�Ћ���E�P���   �	�у�4�M������_^��]������������U������4�@��p  �Ѕ�u��]�Vh#���M��4������M��uh#���@�@4�С���M�j Q�M��@hicMCQ��X  �Ћ�����E�    �E�    j ���   �M�RQ�@�С���M�Q���   � �С���M�Q���   �@8�Ћ�����E�P���   �	�у�(�M���
����^��]�������U������4�@��p  �Ѕ�u��]�Vhs���M��T
������M��uhs���@�@4�С���M�j Q�M��@hicMCQ��X  �Ћ�����E�    �E�    j ���   �M�RQ�@�С���M�Q���   � �С���M�Q���   �@8�Ћ�����E�P���   �	�у�(�M���	����^��]�������U�����@���  ]��������������U�����@���  ]��������������U�����@��@  ]��������������U��V�u���t���Q�@��D  �Ѓ��    ^]�������U�����@��H  ]��������������U�����@��L  ]��������������U�����@��P  ]��������������U�����@��T  ]��������������U�����@��X  ]��������������U�����@��\  ]�������������̡���@��d  ��U�����@��h  ]��������������U�����@��l  ]��������������U�����@���  ]�������������̡���@���  ��U�����@���  ]�������������̡���@��P  �����@���  ��U�����M���@�uQ���  �ЋM��P����M�����E��]���������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@��l  ]��������������U�����@���  ]��������������U�����@���  ]��������������U�����@��$  ]��������������U�����@��(  ]��������������U�����@��,  ]�������������̡���@��0  �����@��<  ��U�����@��  ]��������������U�����@��`  ]��������������U�����@��\  ]��������������U�����u�u�@TQ�@�Ѓ�]� ��U�����uQ�@T�@�Ѓ�]� �����U�����uQ�@T�@�Ѓ�]� �����U�������u�@TQ�M�Q�@<�ЋM���o ��~@��f�A��]� �����U�����@T� ]��U����V�u�@@�6�@�Ѓ��    ^]��������������̡��hG  �@T� �Ѓ�������������U����V�u�@@�6�@�Ѓ��    ^]���������������U�������E�@H�$Q�@�Ѓ�]� ����������̡��j Q�@H���   �Ѓ�����������U�����uj �@HQ���   �Ѓ�]� ���jQ�@H���   �Ѓ�����������U�����uj�@HQ���   �Ѓ�]� ���jQ�@H���   �Ѓ����������U�����uj�@HQ���   �Ѓ�]� ���Q�@H���  �Ѓ�������������U�����uQ�@H���  �Ѓ�]� ��U�����uQ�@H���  �Ѓ�]� ��U�����uQ�@H���  �Ѓ�]� ��U�����u�u�@HQ��  �Ѓ�]� ���������������U�����u�u�@HQ��  �Ѓ�]� ��������������̡��Q�@H���   �Ѓ�������������U��VW�u����  ������t����uV�AHW���   �Ѓ���_^]� �������U��VW�u���u�n�  ������t����uV�AHW���   �Ѓ���_^]� ����U�����u�u�@HQ���   �Ѓ�]� ���������������U�����u�u�@HQ���   �Ѓ�]� ���������������U�����uQ�@H���   �Ѓ�]� �̡��Q�@H���  �Ѓ�������������U���u����u�u�@H�u�u���  Q�Ѓ�]� ������U�������@HWj �����   h�  W�Ѓ��} u�   _��]� Vh�  �_�  ��������   ���j VW�IH���   �у��M��R ������M��uh�  �@�@0�С���M��E���@�$h�  �@,�С���M�j QV�@@�@(�Ѓ��M��Y ��^�   _��]� ^3�_��]� �̡��Q�@H���   ��Y��������������U�����uQ�@H���  �Ѓ�]� ��U�����uQ�@H���  �Ѓ�]� �̡��Q�@H��4  �Ѓ�������������U�����@H� ]��U����V�u�@@�6�@�Ѓ��    ^]���������������U��S�]V�uW�; ���
  ����uW�@H���   �Ѓ�����   ���jW�@H���   �Ѓ�����   ����W�@H���   �Ѓ��} u!�u���S�u�@HV�u���  W�Ѓ��>��t:�u���S�u�@HV�u���  W�С�����΋��   �@(�Ћ���uɋu�; uS���W�@H���   �Ѓ���t;�    ���W�@H���   �С���uW�@H���   �Ѓ�_^[]� �   �   ���W�@H���   �С�����} �@Hu!�u���  j �uV�uW�Ѓ���_^[]� � h  �Ћ؃���u_^[]� ����΋��   �@x�Ћ��P���   �ˋB|�Ѕ�tP�u���j �u�@HV�u���  W�Ћȃ���t���S���   �@H�С���΋��   �@(�Ћ���u�_^��[]� ����U���u����u�u�@H�u�u���  Q�Ѓ�]� �����̡��Q�@H���   ��Y�������������̡��Q�@H���   �Ѓ�������������U�����u�u�@HQ���   �Ѓ�]� ��������������̡��Q�@H���   ��Y�������������̡��Q�@H��t  ��Y�������������̡��Q�@H��P  �Ѓ������������̡��Q�@H��T  �Ѓ������������̡��Q�@H��X  �Ѓ�������������U�������@HQ�M�Q��\  �ЋM���o ��~@��f�A��]� ����̡��Q�@H��`  �Ѓ�������������U�����uQ�@H��d  �Ѓ�]� ��U�������E�@H�$Q��h  �Ѓ�]� ��������U�������E�@H�$Q��t  �Ѓ�]� ��������U�������E�@H�$Q��l  �Ѓ�]� ��������U�����uQ�@H��p  �Ѓ�]� ��U���u����u�u�@H�uQ���  �Ѓ�]� ���������U���u����u�u�@H�u�u���  �uQ�Ѓ�]� ��̡��h�  �@H� �Ѓ�������������U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@H���   �Ѓ������������̡��Q�@H���   �Ѓ�������������U�����uQ�@H���   �Ѓ�]� ��U�����uQ�@H���   �Ѓ�]� ��U�����u�u�@HQ��   �Ѓ�]� ���������������U�����u�E���@H�$���  Q�Ѓ�]� �����U����Vh  �@H� �Ћ�������   �uh�  葆  �Ѓ���t^���j RV�AH���   ���uh(  �f�  �Ѓ���t3���j RV�AH���   �С�����΋��   j j�@�Ћ�^]á��V�@@�@�Ѓ�3�^]�����U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@H��  �Ѓ������������̡��Q�@H��  �Ѓ������������̡��Q�@H���  �Ѓ������������̡��Q�@H���  �Ѓ������������̡��Q�@H���  �Ѓ�������������U�����u�u�@HQ��  �Ѓ�]� ���������������U�����u�u�@H�uQ��   �Ѓ�]� ������������U���u����u�u�@H�uQ��|  �Ѓ�]� ���������U��EV���u����@H���  �'��u����@H���  ���u(����@H���  V�Ѓ���tP�u���   ^]� 3�^]� ����������U���SW����  �؅���   �} ��   ���Vj h�  �AHW��p  �Ћ����h�  W�u�IH���   �������E����   �u3��Ή}��'  ����   �E���P�E�P�u�W��  ��t\�u�;u�T������u�U����ɋD�;D�t-����Hl����P�E�p�A�Ѓ��D����tP����  F;u�~��}��MG�}��  �u;��v���^_��[��]� _3�[��]� U������Vj ��@Hh�  V�u�p  �Ѓ��E���u^��]� �EW��u����@H���  �+��u����@H���  ����T  ����@H���  V�Ћ������6  S���o  ���3�h�  V�]��@H���   �Ѓ�����   �E��s���E����MS�@l�q�@�Ћ؃�����   ����s�u�I\�I,�у���t�F���P�  ����s�u�@\�@,�Ѓ���t�F���P�q  �M�;At"����s�u�@\�@,�Ѓ���tV���E  ����s�u�@\�@,�Ѓ���t�F��P�   ������]��ECh�  �@H�u�]����   �Ѓ�;�����[_�   ^��]� _3�^��]� ������̡��Q�@H���  �Ѓ�������������U�����u�u�@HQ���  �Ѓ�]� ���������������U�����u�u�@H�uQ���  �Ѓ�]� �����������̡��Q�@H���  �Ѓ������������̡��Q�@H���  �Ѓ�������������U�����uQ�@H��  �Ѓ�]� ��U�����uQ�@H��  �Ѓ�]� �̡��Q�@H��  �Ѓ�������������U�����uQ�@H��  �Ѓ�]� �̡��Q�@H��T  �Ѓ�������������U�����u�u�@HQ��  �Ѓ�]� ���������������U�����uQ�@H��8  �Ѓ�]� ��U�����uQ�@H��<  �Ѓ�]� ��U�����u�u�@H�uQ��@  �Ѓ�]� ������������U�����uQ�@H���  �Ѓ�]� ��U�����uQ�@H��H  �Ѓ�]� �̡��Q�@H��L  ��Y��������������U����Vh�  �@H� �Ћ�����u^]á���u�u�@HV��  �Ѓ���u���V�@@�@�Ѓ�3���^]����������U����V�u�@@�6�@�Ѓ��    ^]���������������U�����u�u�@H�uQ��   �Ѓ�]� ������������U�������E�@H�$Q��$  �Ѓ�]� �������̡��Q�@H��(  �Ѓ�������������U�����u�u�@HQ��,  �Ѓ�]� ��������������̡���@H��  ��U�����@H��  ]�������������̡��V��W�@@V�@,�Ћ�����ȋBj h�  ���   �Ћ����h�  V�IH���   �у���
��t_3�^Ë�_^�̡��Q�@@�@,�Ћ�����ЋA��j h�  ���   �����U�������E�u�@H�u����  �$Q�M�Q�ЋM���o ��~@��f�A��]� ��U�������E�u�@H�u����  �$Q�M�Q�ЋM���o ��~@��f�A��]� �̡��Q�@H���  �Ѓ�������������U�����u�u�@HQ��8  �Ѓ�]� ���������������U���u����E���@H�$�u��0  Q�Ѓ�]� ��U�����@H�@]�����������������U����V�u�@@�6�@�Ѓ��    ^]���������������U���u ����u�E���@H�$�u���   �u�u�Ѓ�]�������������U���u����E���@H�$�u�u���   �u�Ѓ�]�����������������    ���������̡��j�1�@H��|  �Ѓ����������U����V�u��@H��x  ��3ɉ��������^]� ���̡��j �1�@H��|  �Ѓ����������U��fnE�M����YE�X���,�;�}��]�;EOE]����������������U���D���SVW�@H�}h�  W���   �Ћ��3�V��h�  �IHW�]ԋ��   �у��E��u��u�u����t	  ����ϋ��   �@��=�  �����  �@HVh:  W���   �Ћ��h�  W�E�IH���   �ы��Vh�  W�IH�E�u؋��   �ы����W�]�IH��  �ы��W�EЋIH���  �у�(�E�3��E�\�9u���   �C3ۉE��MЅ�tNj�W�!�  ���t>�M̍@�|� ���M�~�� ��%�������;�u+蟛  �M�;�O��b�  ���E��M�� ;Au������E�G���E�;}�|��]؋]�E�}����   j W���l~  ���5  �M��~  ��tk�M�� x  �M�;�u\����Ih`���h�  �@Q�Mȋ��  �Ѓ��EĉE�����  �M���}  �Ѕ�t�Eą�t�Mȅ�tQRP�`�  ���E�h`�h�  �@�����Q�Mċ@���  �Ѓ��E����  �U���t�Mą�tQRP��  ���M؅�~,���h`���h�  �@Q���   �Ѓ��E����=  ���j�VW�@H��  �Ѓ����  �u��t jW���<}  ���  ���}  ���E��3��u���j h�  W�@H���   �ЉE�3�3��U����E�9E���  �{�}����$    ��MЅ��  j�P���  ����  �M̍@�|� �4��u�~�� ��%�������9E��2  ���@�  3ۉE�3��E�    9^�{   ��������Шte�E��������������u����E��T��E��N�L��J�E��L��E��N�L��J�E��L��E��N�uȉL��J�E��L���C;^|�����  �ǍM��+�j��P�u�聁  �U�3��]��M��R�ÉE��+ÉEȋƍd$ ;E���  �E�����t.�E��[�oȋM�E���E��[�~D��E�M�f�D�E�[�oȋM���[�~D��M�f�A;�}j�E�9�u_�L�������������w>�$����M���U����-�M���U��T���M���U��T���M���U��T���U���;�|��M�E܃�B�M�M�@�U��E�;�����;E���  �}��_  �U��3�;G�M��Å���   �R�ƋG��@�o���~D�f�B�G��@�E��o��B�~D�f�B(��U��@�E��ȍR�o�D�0�~Af�D�@��t%�G�@�E��oȍȍR�D�H�~Af�D�X�G��u��@�E��oȍȍR���~Af�D��G��W�B�@�E��oȍȍR���~Af�D���W�B�@�E��oȍȍR���~Af�D��B�U���t-�G�@�E��oȍȍR���~Af�D��WB�U����G��}ԋU��E؃��u�@�E؉}�;E��i����E�P�`����E�P�W�������  �E�P�F����E�P�=����E�P�4�����3�_^[��]Ë��   �ϋ@��=  ��  ���j h(  W�@H���   �Ћ����h(  W�IH���   �у��E�3Ʌ�~�I �˅�t�|� �4Vu���A;�|�E�h`�hK  �@�����Q�M��@���  �Ћȃ��M����   �U���t�E���tPRQ躾  ���E�h`�hP  ��    ���Q�M��@���  �Ћȃ��M��tP��t�E���tPSQ�p�  ������ƙ+����IHPVW��   �E��у���u�E�P�����E�P������_^3�[��]á��j h�  W�@H���   �Ћ��j h(  W�IH�E����   �ы�3��E�3ۃ��M�3҉uĉ]܅���   �}�d$ �߅���   3��Eԃ�~d�M��X�R�4v�����E�I0�EԍvC���oD��A��~D�f�A��E��o�A��~D�E�f�A��}�;ǋE�|��uċ]܃|� tL�}�ƍ@�E��oȍȍRB���~A�vf�D��E��oȍȍRB���~Af�D��}�4ߋE؉u�C�]�;������M��U�3���~�I �D�    ��   @;�|�E�P�s������E�P�g�����_^�   [��]�����	����������U���u����E���@H�$�u�u���  �Ѓ�]���U�����@H���  ]��������������U�����@H���  ]��������������U���u0�E(������@H�$�u$�u ���  �u�u�u�u�u�u�Ѓ�,]�U�����@H���  ]��������������U�����@H���  ]��������������U���u0�E�u,����u(�u$�@H�u ����P  �D$�E�$�u�u�Ѓ�,]�������������P����A    ��q�P�����@l�@��Y���������U����V��@l�v�@�ЋM����u�A^]� ����u�u�@lQ�u� ��3ɉF��������^]� �������������̋I��u3�á��Q�@l�@�Ѓ������U�������U�R�U�R�u�@l�u�q�@�ЋM����U;�u	�E���]� ���9U�D���]� �������U�����@H���   ]��������������U�����@H���  ]��������������U���������MW��@�$�u���   ���E�]��M�f/�w�Ef/�w(�������M�@�$�u�@,�Ћ�]����������U���H����M�W�Q�ufE�M��E��@Q�M���   ���M�o �~`�E��Ef/�v(��	f/�v(��U�f/�v(��	f/�v(��]�f/�wf/�v(��(á���M��E��U��e��@Q�u�M�@H�Ћ�]��������U�����@H��0  ]�������������̋������������������������������̡���@H���  ��U�����@H���  ]��������������U���u0����u,�u(�@H�u$�u ���  �u�u�u�u�u�uQ�Ѓ�0]�, ����U���u0����u,�u(�@H�u$�u ���  �u�u�u�u�u�uQ�Ѓ�0]�, ���̡��Q�@H��,  �Ѓ�������������U�����uQ�@H��X  �Ѓ�]� �̡��Q�@H��\  �Ѓ�������������U����Q�u�@H�u���   �Ѓ�]� ���������������U��V���v�P�����@l�@�Ѓ��Et	V�e�������^]� �����������U��E�M� +]� ��������������̡��Q�@\�@�Ѓ���������������̡��Q�@\�@�Ѓ����������������U�����uQ�@\�@�Ѓ�]� �����U�����u�u�@\Q�@�Ѓ�]� ��U�����uQ�@\�@�Ѓ�]� ����̡��Q�@\�@�Ѓ����������������U�����uQ�@\�@ �Ѓ�]� �����U�����u�u�@\Q�@$�Ѓ�]� ��U���u����u�u�@\�uQ�@`�Ѓ�]� ������������U�����uQ�@\�@0�Ѓ�]� �����U�����uQ�@\�@@�Ѓ�]� �����U�����uQ�@\�@D�Ѓ�]� �����U�����uQ�@\�@H�Ѓ�]� ����̡��Q�@\�@4�Ѓ����������������U�����u�u�@\Q�@8�Ѓ�]� ��U�����uQ�@\�@<�Ѓ�]� �����U���SVW�}��j �ω]��������S�@\�@�Ѓ��؋�S����3���~?��I ����M�Q�MQ�@\h���V�u��@`�Ѓ����u�U����u����K���F;�|�_^[��]� �������������U���S�]�E�W����P�����}� |z���W�@\�@�Ѓ��E���P�����E���tWV3���~B�E��P�m����E���P�b����M;M����QW�@\�@�ЋM��A�M;M�~�F;u�|�^_�   [��]� _�   [��]� ����������̡���@\� ������U����V�u�@\�6�@�Ѓ��    ^]��������������̸   � ��������3�� �����������3�� ����������̸   @� ��������3�� ����������̸   � ��������U�����u�H�I�ыE��]� ��̸   � ��������U����   V�u��u3�^��]�h�   ��@���j P��  �E�E��E�E��Eh�   ��@�����@���P�u��`����uǅD��� �j�E�c��E����E�r��E�|��E�w��E�m��E�h��E��������� ^��]��������U����   h�   ��@���j P�d�  �Eh�   �E���@���P�uǅ`���    �uj蛹���� ��]�����U���   SV�u(3�W3��]����w  ����M�@�@<�Ѕ��F  �����E�����   �EP�M�螳������M�Q�@�@�С���M�Wj�hp��@Q�@�Ѓ��E�M�P�e����u��E�Wj�P�E�P��\���P�_?�������P��x���P蘷����P�E�P苷������P�����E���t�E� �� t�M����胳����t��x�������p�����t��\�������]�����t�M̃���M�����t����M�Q����@�@�Ѓ���t�M��$����}� t�u(�u$�u��u�u�u���������E�P�i������V�u$j �u�u�u�p�����������EP�I�I�у���_^[��]Ë�`��`��`��`��`��` ���������������U��M�EQj�u��E�A�������]���������������̸   �����������U��V�u��t���u6j�u���������u3�^]Ë��R����ȅ�t��t��E3�;AOʋ�^]�������V������F    ����@4���   �ЉF��^����������V���v�������@4���   �Ѓ��F    �F    ^��� �������������U����u��U��u�E�    �u�E�    �u�uR�U�R�P�E�3Ɂ}�gnolE���]� �����������U���u����u�u�@4�u�u���   �u�q�Ѓ�]� ̡���q�@4���   ��Y�����������̡���q�@4���   ��Y������������U�����u�q�@4���   �Ѓ�]� ����q�@4���   �Ѓ�����������U���u����u�u�@4�q���   �Ѓ�]� ����������U���u����u�u�@4�q���   �Ѓ�]� ����������U��EQh���u�P���R�q�@4���   �Ѓ�]� ���U�����u�u�@4�q���   �Ѓ�]� �������������V������F    ����@4���   �Ћ�����V���R�A4���   �С�����@4���   �ЉF��^����������V���v�������@4���   �Ѓ��F    �F    ^��U�����u�u�@4�q���   �Ѓ�]� �������������U�����u�u�@4�q���   �Ѓ�]� �������������U�����u�u�@4�q���   �Ѓ�]� ������������̡���q�@4���   �Ѓ�����������U���u����u�u�@4�q���   �Ѓ�]� ����������U�����u�q�@4���   �Ѓ�]� U�����u�q�@4���   �Ѓ�]� U�����u�q�@4���   �Ѓ�]� U�����u�q�@4���   �Ѓ�]� U�����u�u�@4�q���   �Ѓ�]� �������������� �������������U�����u�u�@4�q���   �Ѓ�]� �������������U��M��t�u$��u �u�u�u�u�u�P]�����������U��V���v�������@4���   �Ѓ��F    �E�F    t	V褢������^]� �����������    ���A    �A    �A    ���V��~ u=���t���Q�@<�@�Ѓ��    W�~��t��蛬��W�5������F    _^���������U����E�VP���n�������P�   �M���Y�����^��]���U��V��~ u4h��j;h�j��������t�u�������3��F��u^]� �~ t3�9^��]� ����u�@<� �Ћ��F   ���3�����^]� �����V���F   ����@<�@��3ɉ��^�����������������U��	�����u	�@� ]� �@<�uQ�@�Ѓ�]� �����̃y t�   ËQ��u3�á��R�1�@<�@�Ѓ��������V��~ u=���t���Q�@<�@�Ѓ��    W�~��t������W襠�����F    _^���������U��x������u�@� ]Ë@<�uQ�@�Ѓ�]�������U��x���$V��u����A�0�����uQ�@<�@�Ћ�������I�E�SP�I�ѡ���M�QV�@�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M��� �@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С������[t(�H�uV�I�ы���E�P�I�I�у���^��]Ë@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���uV�@�@�С��V�H�E�P�I�ы���E�P�I�I�у���^��]������������U��x���$SV��u����A�0�����uQ�@<�@�Ћ�������I�E�P�I�ѡ���M�QV�@�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M��� �@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С������t)�H�uV�I�ы���E�P�I�I�у���^[��]Ë@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M����@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С�������?����@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���uV�@�@�С��V�H�E�P�I�ы���E�P�I�I�у���^[��]���U��x���$SV��u����A�0�����uQ�@<�@�Ћ�������I�E�P�I�ѡ���M�QV�@�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M��� �@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С������t)�H�uV�I�ы���E�P�I�I�у���^[��]Ë@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M����@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С�������?����@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M����@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С������������@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���uV�@�@�С��V�H�E�P�I�ы���E�P�I�I�у���^[��]�����������U��x���$SV��u����A�0�����uQ�@<�@�Ћ�������I�E�P�I�ѡ���M�QV�@�@�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M��� �@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С������t)�H�uV�I�ы���E�P�I�I�у���^[��]Ë@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M����@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С�������?����@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M����@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С������������@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���M�Q�@�@�С���M�j j�h��@Q�@�С���M����@j Q�M܋@@Q�M��Ѕ��Mܡ��Q�Ë@�@�С�����������@�M�j�u��@H�С���M�j�j��u�@�u��@L�С���uV�@�@�С��V�H�E�P�I�ы���E�P�I�I�у���^[��]���U��E���x�EȉM]�  ������U�����@<�@]�����������������U��E����u��]�VP�M�赝���E�E�    P�E��E    P�M���������   �u�E���tA��t<��uX����u���   �@H�Ћ���Ѓ��A��V�@x�Ѕ�u+�   ^��]á���u���   �@T��VP�Y�������uՍEP�E�P�M��b�����u�3�^��]��������U���DS3ۍM܉]����VQ�@�@�С���M�Sj�h��@Q�@�С���M�Q�@<�@�Ћ�����E�P�I�I�у���u^3�[��]�WV�M�3�艜���E�P�E�P�M��ɜ�����  ��}���   ����u����   �@T�Ћ�������   ������A�M�Q�@�С���M̃��@Qj�M����   Q���Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M܃��@�u�@x���E���t�E� ��t����M�Q����@�@�Ѓ���t����M�Q����@�@�Ѓ��}� u!�E�P�E�P�M�躛�����������_^[��]Ë}���_^[��]��������������U���@SV�u3ۉ]���u^����M�Q�@�@�С���M�Vj�h��@Q�@�С���M�Q�@<�@�Ћ�����E�P�I�I�у���u^3�[��]�V�M��Ś���E�P�E�P�M�������t�W�}�E�����   ����u����   �@T�Ћ�������   ������A�M�Q�@�С���MЃ��@Qj�M����   Q���Ћ�����E�P�I�I�ы���A�M�QV�@�С���M�Q�@�@�С���M����@W�@x���E��t�E ��t����M�Q����@�@�Ѓ���t����M�Q����@�@�Ѓ��} tA�E�_^[��]Ã�u2�M���t+���Q���   �@H�Ћ���Ѓ��A��W�@x�Ѕ�t��E�P�E�P�M�趙���������_^[��]�������̡���@<�@����̃=�� uK�x���t���Q�@<�@�Ѓ��x�    V�5����t��谜��V�J��������    ^������������3�� �����������3�� �����������3��  ����������̸   � ��������3�� �����������3�� ���������������������������3�� �����������3�� ������������ �������������3�� �����������U���   ������h   j P脟  �u �������u�u�u�uP�)   h   ������P�u�uj
谠����8��]����������U��V�u�u�uj �u�uV������E�����   ǆ�   �ǆ�   ǆ�   8ǆ�   Gǆ�   Lǆ�   Qǆ�   Vǆ�    ǆ�   
ǆ�   =ǆ�   B^]Ë�`P��`X��`\��``��`d��`h��`l����̸   � ��������3�� �����������3�� ������������ �������������U��EW� �@]� �����������3�� �����������3�� ������������ �������������� �������������U������   �M�@�@<�Ѕ�tj �u�u�6�������u��]�h   ������j P蘝  �u �������u�u�uP�    h   ������P�u�uj�Ǟ����4��]�U��V�u�u�uj �u�uV�������ǆ�   �ǆ�    ǆ�   ǆ�   8ǆ�   
ǆ�   =ǆ�   Bǆ�   Gǆ�   L^]Ë�`D��`H��`L��`T�U��Vj j�u����������t�@��t	����^]� 3�^]� U��Vj j�u���~�������t�@��t	����^]� 3�^]� U��Vj j�u���N�������t�@��t����^]� �������U��Vj j�u����������t�@��t	����^]� 3�^]� U��Vj j�u�����������t�@��t	����^]� 3�^]� U��Vj j�u����������t�@��t	����^]� 3�^]� U��Vj j �u����������t�@ ��t�u����^]� 3�^]� �������������U���(Vj j$�u���K�������t^�@$��tW�M�Q���Ћu�Vj �����    �B    ���PR���   �I�ы���E�P���   �	�у���^��]� ����M��E�    �E�    �E������E�    �E�    ���   j Q�M��@Q�С���M�Q���   � �Ћu�E؍Vj ��    �B    ������   �E�PR�I�ы���E�P���   �	�у� ��^��]� �������U��Vj j(�u���.�������t�@(��t�u����^]� ����U��Vj j,�u�����������t�@,��t	����^]� 3�^]� U��Vj j0�u�����������t�@0��t	����^]� 3�^]� U��E�@���@��@���@���@���@���@ ��@$���@(�@,8�@0��@4
]�����3�� ��`0��`<�U��EVW�9�0;�t_3�^]� �P��u ��u9pu9qu��u�9yu�_�B^]� S�Y��u"��u9yu��u3��u/9pu*[_�   ^]� ��t��t;�u�P��t�A��t�;�t�[_3�^]� U���u�e������@]� ������������Vh��j\hD ���|�������t�@\��tV�Ѓ���^�����U��Vh��j\hD ���I�������t2�@\��t+V��h��jxhD �'�������t�@x��t	V�u�Ѓ���^]� ���������U���Vh��j\hD �����������tG�@\��t@V�ЋEh��jdhD �E��E�    �E�    ��������t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��j\hD ���i�������t2�@\��t+V��h��jdhD �G�������t�@d��t	�uV�Ѓ���^]� ���������U��Vh��j\hD ���	�������tZ�@\��tSV��h��jdhD ���������t�@d��t	�uV�Ѓ�h��jhhD ��������t�@h��t	�uV�Ѓ���^]� �U��Vh��j\hD ������������   �@\��t{V��h��jdhD �c�������t�@d��t	�uV�Ѓ�h��jhhD �;�������t�@h��t	�uV�Ѓ�h��jhhD ��������t�@h��t	�uV�Ѓ���^]� �����Vh��j`hD �����������t�@`��tV�Ѓ�^�������U��Vh��jdhD ����������t�@d��t	�uV�Ѓ�^]� �������������U��Vh��jhhD ���i�������t�@h��t	�uV�Ѓ�^]� �������������Vh��jlhD ���,�������t�@l��tV�Ѓ�^�������U��Vh��jphD �����������t�@p��t�uV�Ѓ�^]� ���^]� ���U��Vh��jxhD ����������t�@x��t	V�u�Ѓ���^]� �����������U��Vh��j|hD ���y�������t�@|��tV�u�Ѓ�^]� 3�^]� ������U��Vh��j|hD ���9�������t�@|��tV�u�Ѓ����@^]� �   ^]� ��������������U���Vh��jthD �����������tP�@t��tI�u�M�VQ�Ћu����P�`���h��j`hD ��������th�H`��ta�E�P�у���^��]� h��j\hD �~����u����t4�@\��t-V��h��jdhD �Y�������t�@d��th��V�Ѓ���^��]� �������U��Vh��h�   hD ����������t���   ��t�uV�Ѓ�^]� 3�^]� U��Vh��h�   hD �����������t���   ��t�uV�Ѓ�^]� 3�^]� VW��3����$    �h��jphD ��������t�@p��t	VW�Ѓ������8 tF��_��^�������U��SV��3�W��    h��jphD �?�������t�@p��t	VS�Ѓ������8 tph��jphD ��������t�@p��tV�u�Ѓ�������h��jphD ���������t�@p��t	VS�Ѓ�����W���x�����tF�^����E_��t�0��~=h��jphD ��������t�@p��t	VS�Ѓ������8 u^�   []� ^3�[]� �����������U���Vh��h�   hD ���3�������t<���   ��t2�u�M�VQ��h��j`hD ��������t�@`��t	�M�Q�Ѓ���^��]� �������U���Vh��h�   hD ���������tS���   ��tI�u�M��uQ�Ћu����P�:���h��j`hD ��������td�H`��t]�E�P�у���^��]�h��j\hD �Z����u����t2�@\��t+V��h��jxhD �5�������t�@x��t	V�u�Ѓ���^��]�������̋���������������h��jhD ���������t	�@��t��3��������������U��V�u�> t+h��jhD ��������t�@��tV�Ѓ��    ^]�������U��} W��t0h��jhD �s�������t�@��t�u�uW�Ѓ�_]� 3�_]� �������������U��Vh��jhD ���)�������t�@��t�uV�Ѓ�^]� 3�^]� ������U��Vh��jhD �����������t�@��t�uV�Ѓ�^]� 3�^]� ������Vh��j hD ����������t�@ ��tV�Ѓ�^�3�^���Vh��j$hD ���|�������t�@$��tV�Ѓ�^�3�^���U��Vh��j(hD ���I�������t�@(��t�u�u�uV�Ѓ�^]� 3�^]� U��Vh��j,hD ���	�������t�@,��t�u�uV�Ѓ�^]� 3�^]� ���U��Vh��j(hD �����������t�@0��t�u�u�uV�Ѓ�^]� 3�^]� Vh��j4hD ����������t�@4��tV�Ѓ�^�3�^���U��Vh��j8hD ���Y�������t�@8��t�u�u�u�uV�Ѓ�^]� 3�^]� �������������U��Vh��j<hD ���	�������t�@<��t	�uV�Ѓ�^]� �������������U��Vh��h�   hD �����������u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ����������u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ���F�������u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ����������t�u���   �u�uV�Ѓ�^]� �����Vh��jDhD �����������t�@D��tV�Ѓ�^�3�^���U��Vh��jHhD ����������t�u�@HV�Ѓ�^]� �U��Vh��jLhD ���i�������u^]� �u�@LV�Ѓ�^]� ������������U��Vh��jPhD ���)�������u^]� �u�@P�uV�Ѓ�^]� ���������U��Vh��h�   hD �����������u^]� �u���   �u�uV�Ѓ�^]� U��Vh��h�   hD ����������u^]� �u���   �u�u�u�uV�Ѓ�^]� ����������Vh��jThD ���\�������u^Ë@TV�Ѓ�^���������U��Vh��jXhD ���)�������t�u�@XV�Ѓ�^]� �U���Vh��h�   hD �����������tQ���   ��tG�u�M�Q���Ћu��P�l���h��j`hD ��������t|�H`��tu�E�P�у���^��]� h��j\hD �E�    �E�    �E�    �u����u����t3�@\��t,V��h��jdhD �P�������t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��h�   hD ����������t���   ��t�u���u�u��^]� 3�^]� ������������U��Vh��h�   hD ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   hD ���v�������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   hD ���6�������t���   ��t�u����^]� 3�^]� ��Vh��h�   hD �����������t���   ��t��^��3�^����������������U��Vh��h�   hD ����������t���   ��t�u���u�u��^]� 3�^]� ������������U��Vh��h�   hD ���f�������t���   ��t�u����^]� ���������U��Vh��h�   hD ���&�������t���   ��t�u���u�u��^]� 3�^]� ������������Vh��h�   hD �����������t���   ��t��^��3�^����������������U��h��jhD ��������t
�@��t]��3�]��������U���Vh��h�   hD �e�������u����uV�H�I�у���^��]Ë��   �M�W�uQ�Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]���U��h���uhD �������]�������Vh��h�   h D ����������t���   ��t��^��3�^����������������Vh��h�   h D ���y�������t���   ��t��^��3�^����������������Vh��h�   h D ���9�������t���   ��t��^��^��U��Vh��h�   h D ����������t���   ��t�u����^]� 3�^]� ��Vh��h�   h D �����������t���   ��t��^��^��U���Vh��h�   h D ����������t=���   ��t3�E�M���$Q���ЋM^�o ��~@��f�A��]� �EW�^ �@��]� ����������Vh��h�   h D ����������t���   ��t��^��3�^����������������U��Vh��h�   h D �����������t���   ��t�u����^]� ���^]� �U��Vh��h�   h D ����������t���   ��t�u����^]� 3�^]� ��U���8Vh��h�   h D ���S�������tG���   ��t=�u�M�Q���ЋM^�o ��o@�A�o@ �A �~@0��f�A0��]� �EW�(����^�@0    � ���f�H�H�P �@(��]� ���������������U��Vh��h�   h D ����������t���   ��t
�u���u��^]� ������U���Vh��h�   h D ���S�������tZ���   ��tP�u�M�Q���Ћuj PV�    �F    ������   �I�ы���E�P���   �	�у���^��]� �E^�     �@    ��]� �����������U��Vh��h�   h D ����������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h D ���f�������t���   ��t�u����^]� 3�^]� ��Vh��h�   h D ���)�������t���   ��t��^��3�^����������������Vh��h�   h D �����������t���   ��t��^��3�^����������������Vh��h�   h D ����������t���   ��t��^��3�^����������������Vh��h�   h D ���i�������t���   ��t��^��3�^����������������Vh��h�   h D ���)�������t���   ��t��^��^��U��MVh!D �u��������t+h��h�   h D ���������t���   ��t��^]��^]���������h��h�   h D ��������t���   ��t��3��������U��h��h�   h D �y�������t���   ��tV�u�6�Ѓ��    ^]ËE�     ]����������Vh��h�   h D ���)�������t���   ��t��^��3�^����������������U��Vh��h�   h D �����������t���   ��t�u����^]� ���^]� �U��Vh��h�   h D ����������t���   ��t
�u���u��^]� ������U��h���uh D �k�����]�������U��U�f.���D��   �Af.B���D��   �Af.B���Dzy�A;Buq�A f.B ���Dza�A(f.B(���DzQ�A0f.B0���DzA�A8f.B8���Dz1�A@f.B@���Dz!�AHf.BH���Dz�A;Bu	�   ]� 3�]� �����U���u�5������@]� ������������h��h  h�e �l�������t��  ��t��3��������U��h��h  h�e �9�������t��  ��t]��]����Vh��h�   h�e ���	�������t���   ��t��^�����^���������������U��Vh��h�   h�e �����������t���   ��t�u����^]� 3�^]� ��U���Vh��h�   h�e ����������t=���   ��t3�E�M���$Q���ЋM^�o ��~@��f�A��]� �EW�^ �@��]� ����������Vh��h�   h�e ���	�������t���   ��t��^��^��U��Vh��h�   h�e �����������t���   ��t�u����^]� 3�^]� ��U��Vh��h$  h�e ����������t��$  ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ���V�������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e �����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ���V�������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e �����������t���   ��t�u����^]� 3�^]� ��U��Vh��h  h�e ����������t��  ��t�u���u��^]� 3�^]� ���������������Vh��h  h�e ���I�������t��  ��t��^��^��Vh��h�   h�e ����������t���   ��t��^��^��Vh��h�   h�e �����������t���   ��t��^��^��Vh��h�   h�e ����������t���   ��t��^��^��Vh��h�   h�e ����������t���   ��t��^��^��U��Vh��h  h�e ���V�������t��  ��t�u���u��^]� 3�^]� ���������������U��Vh��h   h�e ����������t��   ��t�u���u��^]� 3�^]� ���������������U��Vh��h<  h�e ����������t��<  ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ���v�������t���   ��t�u����^]� ���������Vh��h�   h�e ���9�������t���   ��t��^��3�^����������������U��Vh��h  h�e �����������t%��  ��t�u���u�u�u�u�u��^]� 3�^]� ���U��Vh��h  h�e ����������tR��  ��tH�E0��0���D$(�E(�D$ �E �D$�E�D$�E�D$�E�$��^]�0 ��������U��Vh��h(  h�e ���&�������tR��(  ��tH�E0��0���D$(�E(�D$ �E �D$�E�D$�E�D$�E�$��^]�0 ��������U��Vh��h�   h�e ��覿������t.���   ��t$�u�E�΃��D$�E�$��^]� ���^]� ���������U��Vh��h�   h�e ���F�������t���   ��t�u����^]� 3�^]� ��U��Vh��h0  h�e ����������t��0  ��t�u����^]� 3�^]� ��U��Vh��h,  h�e ���ƾ������t��,  ��t
�u���u��^]� ������U��VWh��h�   h�e ��腾��������tG���    t>j<j h���ut  ����� ;���0;�ϋ��   �uh��j<h����_^]� ���������������Vh��h�   h�e ���	�������t���   ��t��^��3�^����������������U��Vh��h�   h�e ���ƽ������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�e ��膽������t���   ��t�u����^]� ���������U��Vh��h�   h�e ���F�������t���   ��t�u����^]� ���������Vh��h�   h�e ���	�������t���   ��t��^��3�^����������������Vh��h�   h�e ���ɼ������t���   ��t��^��3�^����������������U��Vh��h   h�e ��膼������t ��   ��t�u���u�u�u�u�u��^]� ����������U��Vh��h4  h�e ���6�������t��4  ��t�u���u�u��^]� ���U��Vh��h8  h�e �����������t��8  ��t�u���u�u��^]� ���U��M���E��D$�E�$�]� ����������U��M���E��D$�E�$�u�P]� ������U��h���uh�e �[�����]�������U��h��jhD �<�������t
�@��t]��3�]��������U��h��jhD ��������t
�@��t]��]����������U��h��j8hD �ܺ������t
�@8��t]��]����������U��QVh��j8hD 誺��������th�~8 tb������   ���   �ЉE���t-����u���   �ȋ��   ���u�F8�u�u��u�Ѓ�����M�Q���   ���   �Ѓ�^��]�����h��jhD ��������t	�@��t�����������������U��h��jhD ��������t
�@��t]��3�]��������U��V�u��u3�^]á�����   ���   �ЉE��tF���V���   �ȋ��   �Ћuh��jhD �{�������t�@��t�uV�Ѓ����3�����MQ���   ���   �Ѓ���^]����������������U��h��j4hD ��������t
�@4��t]��3�]��������U��h��j hD ��������t
�@ ��t]��3�]��������U��h��j$hD 輸������t
�@$��t]��3�]��������h��j(hD 菸������t	�@(��t��3��������������U��h��j,hD �\�������t
�@,��t]��3�]��������h��j0hD �/�������t	�@0��t��3��������������U��h���uhD �������]�������h��jhD �߷������t	�@��t��3��������������U��h��jhD 謷������t
�@��t]��3�]��������U���(t��������u�u�A�ʋ��   �ЋE�袅���} tj�r����]� j �wr����]� U��U��3ɋ���tvV�u;�t�D�A���u�^��]� �D����tS�E�   �E��s������ЋA�M�Q�u�ʋ��   �С���M�Q���   � �ЋE�����j ��q����^��]� ��U���Hs��������u�A�ʋ@t�Ћ��j P�u���   �A�ЋE���]� ���������������U���V��r��������u�A�ʋ@t�Ћ��P���   �@8�ЋU����3��:�tZ��9qt@�<����u�^��]� �M��E�����E�   j Q���   �u�@�С���M�Q���   � �ЋE���^��]� �������������U���V�u�E�    W����   �}��u�*r��������E�    �E�    S�A�ϋ]S�@t�Ћ���Ћ��   �M�QR�@�Ѓ���uC�����S�@�@t�Ћ��P���   �@�Ћ�����u���   �I�у�;�u2�������M�Q���   � �Ѓ���[td������u�u�@���   ��_^��]� ���O����}��tj P���N�����t(j W�������Ѕ�t����uj�A�ʋ��   ��_^��]� ����������V���c������^���������������U��V�uj �u�uj �uV��   ����u3�^]�j#V��c��������t���V�@@�@,�Ћ�����ЋA���uh�  �@4�С��V�@@�@,�Ћ�����ЋA���uh�  �@4�Ћ�^]���������������U��h���uhD 蛳����]�������U��V�uW�u�}j W�u�uV�#��������   _^]�������U������   �@V�u�΋@<�Ѕ�tj V�u���������u^��]�h   ������j P�&i  �u������j j V�u�uP謓��h   �������u�P�u�uj#�Pj����8^��]���������Vh��jh�t���輲������t�@��t��^��3�^������Vh��jh�t���茲������t�@��t��^��3�^������U���Vh��jh�t����V�������tV�@��tOW�u�M�Q���Ћ�����}W�I�I�ы��WV�I�I�ы���E�P�I�I�у���_^��]� ����uV�H�I�у���^��]� ������������Vh��jh�t���輱������t�@��t��^��3�^������U��Vh��jh�t���艱������t�@��t�u���u��^]� 3�^]� �����U��Vh��j h�t����I�������t�@ ��t�u���u��^]� 3�^]� �����Vh��jh�t�����������u^Ë@V�Ѓ�^���������U��h���uh�t��۰����]�������U��Vh��h�   h�f ��趰������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h�f ���f�������t���   ��t�u���u��^]� ���^]� ��������������U��Vh��h�   h�f ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�f ���֯������t���   ��t
�u���u��^]� ������U��Vh��h�   h�f ��薯������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�f ���V�������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h�f ����������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h�f ��趮������t���   ��t�u����^]� 3�^]� ��Vh��h�   h�f ���y�������t���   ��t��^��3�^����������������U��Vh��h�   h�f ���6�������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h�f �����������t���   ��t�u���u��^]� 3�^]� ���������������Vh��h�   h�f ��詭������t���   ��t��^��3�^����������������U��Vh��h�   h�f ���f�������t���   ��t�u����^]� 3�^]� ��U��V�u�> t2h��h�   h�f � �������t���   ��t�6�Ѓ��    ^]����������������U��h���uh�f �۬����]�������U��E���� ]��U��EHV����   �$�K�   ^]á �@� �����   �u������=�2  }�����^]Ëu��t�hh�jmh�j�hW������tl���]�������tfV���9b���   ^]��u�u�6����������H^]�^]�a���� �u.������_����5����t���>^��V��S�������    �   ^]Ã��^]Ð0J�J�J(J�J�J����U���Mu�E����E����   ]� ��������������̋ыB�����t!�J��t�H�J�B�A�B    �B    ����������������U��U�B�A�J�A�Q�H]� ����U��U�B�A�J�A�Q�H]� ���̋ыB��t!�J��t�H�J�B�A�B    �B    ����������Q����A�B    �B    � ���@    �@    �A���A    �A    �Q�A    ���������������V������  �N�F����t!�F��t�A�N�F�A�F    �F    �N�F����t!�F��t�A�N�F�A�F    �F    ^���U��A3҃�V;�t��t�u��B;�t�@��t
�x t��u�3�^]� ����������U��U�A�B�A�B�A�P�Q]� �U��U�A�B�A�B�A�P�Q]� ̍A�A    �A�A�A�A    ������SW���O�_;�t!��tV�q��t�~ u3��j��΅�u�^�G�_�G    �G�G    _[�������̋A��;�tE��tAV��H��t
�y t���3��P��t��t�J�P�H�J�@    �@    �ƅ�u�^ËQ�AV3�;�t��t�RF��t
�z t��u��^����������VW���w���V��R�����G    �G    �    _^����U��S�]V��F;�~ ��x�N�E^���   []� ^3�[]� }hW�~9~uI��u�~��F��t�����t?���h��j8�H��    P�v��  �Ѓ���t�F�~�N�F��    �F9^|�_�F;Fu����  ���w����V�N�E���   �F^[]� ����U��UV���x'�F;�} �M��x;�};�t�F���4��
���^]� �������U��UV�uW��;�}N��x.�G;�}'��x#;�};�t�GSR���j  ��t	VS����   [_^]� ������U����Ej�q�E���q�M��E���  ��]� �������U����Ej�q�E���q�M��E��u��  ��]� ����VW���O�q���x6;�}2�G����t*��x&;�}"�w;�}��I �O��F�J�
;w|�_^�3�_^��������U��V��F;Fu�}  ��u^]� �V�N�E���   �F^]� �����������U��V��W�}�F;�O�3Ʌ�H�;Fu���+  ��u_^]� �F;�~�N��H�J��
;���N�E���   �F_^]� ���U��UV���x.�F;�}'H�F;�}�d$ �F��B�A�;V|�   ^]� 3�^]� ��������������U��V��3�W�N��~�V�}9:t@��;�|�����x(;�}$I�N;�}�N��@�J�
;F|�_�   ^]� _3�^]� �������U��Q3�V��~�I�u91t@��;�|���^]� ����������A    ���������VW���wV�#O�����G    �G    �    _^����������U��QSV�uW���}��FP��N���V�F    �    3��F    ���G�F�G�F9_~r�G�~���E9~uJ��u�~��F��t�����tU���h��j8�H��    P�2��  �Ѓ���t-�V�~��NC��}�<��}��F;_|�_^�   [��]� _^3�[��]� V��W�~��u�~��F��t�����u_3�^á��h��j8�H��    P�v��  �Ѓ���t҉~�F�   _^����U��VW���w���V�M�����    �E�G    �G    t	W�K������_^]� ������������U��V�������Et	V��J������^]� ���������������U��V��F�����t!�N��t�H�N�F�A�F    �F    �Et	V�J������^]� ������U���u�A�u�Ѓ�]� �����������U��h�jh�f �\�������t
�@��t]�����]�������U��Vh�jh�f �+���������t=�~ t7�u8�E�u4�u0�u,�u(����P�T���u�F�Ѓ�4�M���:T����^]ÍM����*T����^]������U��h�jh�f 輡������t
�@��t]��3�]��������U��h�jh�f 茡������t�x t�@]��3�]������U��h��uh�f �[�����]�������U������V���.�vf(�fT@�f(�f/�fT@��U��M��M��  f/��  �`�f/�vFf/�v@�,��,���   ��$    ������ʅ�u�fn�����^��^��.�v^��]�f/�v(��(��p��^��%��f/�v1(��Y��Y��Y��.�E�(��Y��v(��M��M�f/�v(��f�E��E���    �E��E��1  �M��]��E�f/��f��M��E��E�s�f^�^��]�W������F^��]����U���E�h�f/�V��w�x�f/�v(��Y�����X���E�E�$�N  ��������F�������^]� ���U����M3��UW�f/�V��fT@��X����3�f/��M��E���3�;������M�$�M  �EfT@��E�X����E�E�$�oM  ������]�Ef/��Fv'���h�j�@��0  ��������F�} u�fWP�����-�����^��]� ����U���E���f/�V���Fv'���h�j,�@��0  ��������F^]� ������U���M�����f/�V��v'���h�j5�@��0  ��������M����Y��E��E��$�RL  �]��F�$�DL  �E��]��^E��E��E��$�'L  ��E�$�L  �����^�-���^��]� �����̡��Q�@D�@$�Ѓ����������������U����j �u�@D� �Ѓ�]��������U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�����@D� ]��U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�����uh2  �@D� �Ѓ�]�����U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@�Ѓ����������������U����j �u�@D� �Ѓ�]��������U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�����uh'  �@D� �Ѓ�]�����U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�����uhO  �@D� �Ѓ�]�����U����V�u�@@�6�@�Ѓ��    ^]���������������U�������@XQ�M�Q� �ЋM���o ��~@��f�A��]� ���������U�������@XQ�M�Q�@�ЋM���o ��~@��f�A��]� ��������U�������@XQ�M�Q�@�ЋM���o ��~@��f�A��]� ��������U������`�@XQ�M�Q�@�ЋM���o ��o@�A�o@ �A �o@0�A0�o@@�A@�o@P���AP��]� U�����uQ�@X�@�Ѓ�]� �����U�����uQ�@X�@�Ѓ�]� �����U�����uQ�@X�@�Ѓ�]� �����U�����uQ�@X�@�Ѓ�]� �����U�����uQ�@X�@$�Ѓ�]� �����U�����uQ�@X�@ �Ѓ�]� ����̡��j h�  �@D� �Ѓ�����������U����V�u�@@�6�@�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�����u�u�@DQ�@�Ѓ�]� �̡��j h:  �@D� �Ѓ�����������U����V�u�@@�6�@�Ѓ��    ^]���������������U�������U��E�    �E�    R���   j�@�����#E���]�����������̡��j h�F �@D� �Ѓ�����������U����V�u�@@�6�@�Ѓ��    ^]���������������U��E����u��]� �E��U�����E�    Rj���   �@������؋�]� ̡��j h�_ �@D� �Ѓ�����������U����V�u�@@�6�@�Ѓ��    ^]���������������U���$�U�M���$  �M�B�S������C�M�VW�}�s��]����Oǉu��]��E��~��}���u��}��~u�K+��]�u��}��9�Ћ��t+��D�R�
��Nu�M�E��UJ�U����   �u�+��E��<�}�;����    �ލw���]�u;�}�U��Q�M���V����y�u�G�}�M�VS���M���U�]�E��Q����F��م�t�}�+���@���T�Ku�}�M�U��}�;�~��]�E�����_^[��]� �U���(SV�u�މM��M���]���8  W����G�}�G���E�E��A����E�����E�E�Ѓ��u�ډU��U��u���}�u���~�u�Ou�)E�}�u��J�֋��t,�}�+}����    f�D�R�
f�f�Nu�M�E�}�I�M����   )E��U��u���}�;���I �ލw����]�u;�}��Q�M܋�V���y�u�G�}�M�VS���M���U��E�]��E����ˍF���t�}�+�f��@�f�f�T�Ku�}�M��U��E�}�;�~��]�����_^[��]� ���������������U���(SV�u�މM��M���]���5  W����G�}�G���E�E��A����E�����E�E�Ѓ��u�ډU��U��u���}�u���~�u�Ou�)E�}�u��E�֋��t'�}�+}���$    �J�R���Nu�M�E�}�I�M����   )E��U��u���}�;����$    �ލw����]�u;�}��Q�M܋�V���y�u�G�}�M�VS���M���U��E�]��F����ˍF���t�}�+��P�@�L���T�Ku�}�M��U��E�}�;�~��]�����_^[��]� �U��U��u	�U]����3������t	�U]�����U]�������������������U��Q�E�M�SW��t*�]��t#�}��t�} t�SP���u
_��[��]� y
_3�[��]� �   O�EV;�|1�M��4�����]�]S�u���ty�E�~���F�E;�~�^_3�[��]� ��~-�M�������؉E}�M��W�uN����u	�E�߅��^_��[��]� ������U����ESVW���}�����   �]����   �u����   �} ��   �SP�����   y�E_^[�     3���]� �N��   3��U�M�;�|6��4���ϋ��]]S�u���t/y�U�N��M��	�M��V�U;�~ʅ��E~F_�03�^[��]� ��~,�E���}�؉E}�M��W�uN����u	�E�߅��_^��[��]� �E_^[� ����3���]� ������    ���A    �A    �A    ���V��V�79���FP�.9�����F    �F    ^������������U��V��W�}j�    �F    �F    �F    �G;Gu2j�   ��tY�����G�A��G_�A�F�    ��^]� j�   ��t'�����G�A��G�A��G�A�F�    _��^]� �����U��V�u���    �F    �F    �F    �  ��^]� U��V�u���  ��^]� �����������U��SV��V�8���FP�
8���]���F    �F    ��t(���h��jI�H��    P���   �Ѓ����u^3�[]� W�}��t;���h��jN�H��    P���   �Ѓ��F��uV�7����3�_^[]� �~�   _�^^[]� �������������V��V�W7���FP�N7�����F    �F    ^������������U��SV��WV�"7���^S�7���}���F    �F    ����   �? ��   �W����   ���h��jl�H��    P���  �Ѓ����t<� t?�W��t8���h��jq�H��    P���  �Ѓ����u���%���_^3�[]� �G��F�G�F�����t��t��tPRQ�;  �����t�FQ��PQ�w�{  ��_^�   []� ������������U��SV��WV�6���~W�	6�����F    �} �F    ��   �]����   �����    h��h�   Q�@���  �Ѓ����t?�} tJ�U��tC���h��h�   �H��    P���  �Ѓ����u������_^3�[]� �E�F�,�F   ���h��h�   j�@���  �Ѓ����t���^��t��    ��tQ�uP�n:  ���U��t ��FQ��PQR�C  ���   _^[]� ��_^�   []� �����    �A    �A    �A    �����U�������   �U��WɉD$VW�H�L$P�L$H�D$    �<��L$}
��_^��]� �u�}���`  �W�f(�f�$�   ��T$(�@�o$��~\��A(�f��d$X�@�\$@���D��\��|��\ŋD$�\�)l$0�f��L$p����   ��$�   ���D$ �����$�   �D$��	��$    ���\$@�f(��L$x���T$p�@�4��\��d��\��l��\�(��Y��Y��Y��Y�f��\�f(��Y��Y��X\$�\��od$X�\��\$�X|$ �t$p�XT$((�f�(l$0�L$ �T$(J�S������$�   ��$�   �L$ �\$W��f�F(��Y�(��Y��X�f(��Y��X���4  �L$W��T$ �|$(f.ş��Dz	W�f(��2����^�f(��Y��D$pf(��Y��Y��D$xfD$p�FHf�^X�@�fT�fT�f/���   f(�fT�f/���   �FH�VX(��fP(��Y��Y��Y��\��\��\�f��^f�f(�~P�NX(��n (��YV(�vH�Y��\�(��YF(�Y��T$0�Vf(��Y��Y��\��   fT�f/��VX��   �FP�NH(��Y��Y��\��\��Y��\�f��^f�N(�f(�n (��YNP(��YFX�vH�\�(��Y��Y��L$0�Nf(��YNP�Y^X�\��\��oD$0f��F0f�v@�   �NPf(��Y�(��Y��\��FH�Y����\��\�f��^0f�F@(��fX�YF@(��YN8�v0�\�(��Y��Y��L$0�NHf(��YN8�Y^@�\��\��oD$0f��Ff�v(��$�   VP�A-���U���o ��o@�F�o@ �F �o@0�F0�o@@�F@�o@P�D$�FP3Ʌ�~w��rr�@�D$��%  �yH���@�T$W�)D$foʋD$���$    ��o�f���oD���f��;L$|�f��fo�fs�f��fo�fs�f��f~L$�D$     �D$    ;�}s��+���|A�D$�@�D$�B��t$�D$ 3�3����$    �|���;L$ |��u�|$�}�D$ ;�}�D$�T$�@��T$�U�D$ D$�L$���L$�D$�F0�V �D$@� �D$�~(�v@(ϋ��@�YD����d�f(��Yn�Y��Y��X.�XV�XN�X��FH�Y��X��F8�YD��X��FP�Y��X�(��YD��D$f�D��X��FX�Yč@�$��\��X��T�(ËD$�l$X�n0f�L$h(��YN�@�Y��X��3��T$�D$ �X�(��YFH�X�(��YF8�Y��L$0(��Y��YN �o|$0�Xf�XN�X��X�(��YFP�YVX�X��X�f�f�d$(���  ���f(��|$�D$ы��@���T�f(��Yv(��\��YŋD$ �X6�n @�Y�D$ �Y�(��X�(��YFH�Xn�Xff��X��F8�Y��X��FP�Y��X��F@�Y��T$`�X��FX�Y�(��\��\��X�f(��\��Y��Y��YD$X�|$X���X�f��l$@�X��X\$P(��D$P�D$H�~D$(f�D$hf�d$(;D$������D$H_^��]� ���U�������������U�   @t������@��wg�$�hu�E� ����E� ���]� �E�
��E�J�]� �E�J��E�J�]� �E�J��E�J�]� �E�J��E�
�]� ��uu+u?uSu����U��S��VW�����%�����   @t�����ʃ��};�t�����t�u�����t��u;�t?�����t7�΁����Eǃ��t����   �_�^�[]� ��   ���Ё�   @�_^[]� �U������4�AW��$W��T$SfD$ V�\$,�L$$�\$�L$W���S  �9�u��$    ������Ш�)  ���������U��Z�@�[�<��l��\<��\l�;Zuc�\��B�\\��@�d��\d��T��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��Xd$(��d�d��B�\d��@�B�@�T��\��\\��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��X\$�XL$�Y��Y��\$�L$�\��Xt$ (��T$ ���L$�����f(��Y�f(��Y��X�f(��Y��X��t+  f(�W�f.П��D�Ez �@_^[��]� ����^�_^[(��YD$� (��YD$�@�D$�Y��@��]� U���<(0��A�=���%��V�E�3��E�(`��E܅��  �m��u��U��E�S��MW��    ������Ш�n  ���������U��@��tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��EċB�@��tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��Eċz���tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��EċB;���   �@��tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��Eă��M��u���_[��ta�Ef(�f(��X�����X�f(��X�^�Y��Y��Y�f��f�P�\0�\h�\`�Ef��0f�`��]� �EW�W�^� f�H�E� f�H��]� ��������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}���x(���t"�v3Ʌ�~�I ���%���;�tA��;�|�_���^]� _��^]� ���������U��SV�q2�3҅�~9W�9����%���;Eu ����   @u�����t	�   ���3�
�B;�|�_��^��[]� ������������V�q3҅�~�	�d$ ��   @u	�����tB��Nu��^�����V�q3҅�~�	�d$ ����ШtB��Nu��^�����������U���V��3�9N~��$����A;N|�N��~kS�   3�W�U��]�����x:�������;�}+�I ����<����������;�u��   ��@;F|ۋU��]�B�N���]��U��B�;�|�_[^��]�����������h�jh_� ��x������uË@����U��V�u�> t/h�jh_� ��x������t��M�M�@Q�Ѓ��    ^]���U��Vh�jh_� ���x������t�@��t�u����^]� 3�^]� ��������U��Vh�jh_� ���Ix������t�@��t�u����^]� 3�^]� ��������U��Vh�jh_� ���	x������t�@��t�u���u�u��^]� 3�^]� ��U��Vh�jh_� ����w������t�@��t�u����^]� 3�^]� ��������U��Vh�j h_� ���w������t�@ ��t�u����^]� 3�^]� ��������U��Vh�j$h_� ���Iw������t�@$��t�u����^]� 2�^]� ��������Vh�j(h_� ���w������t�@(��t��^��3�^������Vh�j,h_� ����v������t�@,��t��^��3�^������U��Vh�j0h_� ���v������t�@0��t�u����^]� 3�^]� ��������U��Vh�j4h_� ���iv������t�@4��t�u���u��^]� ���^]� ����Vh�j8h_� ���,v������t�@8��t��^��3�^������U��Vh�j<h_� ����u������t�@<��t�u����^]� ���������������U��Vh�j@h_� ���u������t�@@��t�u����^]� ���������������U��Vh�jDh_� ���yu������t�@D��t�u����^]� 3�^]� ��������U��Vh�jHh_� ���9u������t�@H��t�u����^]� ���������������Vh�jLh_� ����t������t�@L��t��^��3�^������Vh�jPh_� ����t������t�@P��t��^��3�^������Vh�jTh_� ���t������t�@T��t��^��^��������Vh�jXh_� ���lt������t�@X��t��^��^��������Vh�j\h_� ���<t������t�@\��t��^��^��������U��Vh�j`h_� ���	t������t�@`��t�u���u��^]� 3�^]� �����U��Vh�jdh_� ����s������t�@d��t�u���u��^]� 3�^]� �����U��Vh�jhh_� ���s������t�@h��t�u���u�u�u�u��^]� ���U��Vh�jlh_� ���Is������t�@l��t�u���u�u��^]� 3�^]� ��U��Vh�jph_� ���	s������t�@p��t�u���u��^]� 3�^]� �����U��Vh�jth_� ����r������t�@t��t�u���u��^]� 3�^]� �����U��Vh�jxh_� ���r������t�@x��t�u���u��^]� 3�^]� �����U��Vh�j|h_� ���Ir������t�@|��t�u����^]� 3�^]� ��������U��Vh�h�   h_� ���r������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh�h�   h_� ���q������t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh�h�   h_� ���fq������t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh�h�   h_� ���q������t���   ��t�u���u�u�u��^]� 3�^]� ���������U��Vh�h�   h_� ����p������t���   ��t�u����^]� 3�^]� ��U��Vh�h�   h_� ���p������t���   ��t�u����^]� ���������U��Vh�h�   h_� ���Fp������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh�h�   h_� ����o������t���   ��t�u���u�u��^]� 3�^]� ������������U����M�U�E�A�R�X�\B�\��\Y�Y �Y�Y�X��X��U��E���]�����U��h��uh_� �[o����]�������U��E��t�M��t�U��tRPQ��  ��]��5 �����t��jj �03  YY�H3  U��� SW3ۍ}�j3��]�Y�9Eu�C  �    ��4  ����M�E��t�V�E�E��EPS�u�E��E����P�E�B   �6  �����M�x�M����E�PS�4  YY��^_[��]�;�u���C  �����̺���E  ����D  ���������z�����������������̃=H� t-U�������$�,$�Ã=H� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̃��\$�D$%�  =�  ��  �<$f�$f��f����  f$f%�f fW�f���fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU0fV�f($�0����X��\��Y��Y��Y����X��^�f�f-��\�fs�?��fs�?�Y�fp�Df5��Y��Y�fW��Y�f\%0�Y��X��Y��\�fp���X��\��\ă��-�  ��A�   fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<�0�Y��Y��Y��\�fT@�X��\��X�f-��\��X�f��^�f�fX�0����Y��Y��Y��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fWƃ���;  = 8  ��   f�f(5�f�f(�f(%�fY�f(-0fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��XŃ��-�;  ����   fW�fT=�f%f(��Y�f(��\�f(�fp�D�Q�fY�fp�Df��fY�fX�fpfY�����Y�fX�fp�D�Y�fT@fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^�fX�fY�fp���X�% �  f��fp���X��X��X��X�fWƃ���� = � ��   f~�fs� f~�������  �?+���� ttf$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$��D  fD$�� �f������fn�fp� fPfXfT�fT��X��f0f8�X��fW��Xƺ�  �t���f�$��G  �$�~$��Ð���\$�D$%�  =�  ��  �<$f�$f��f����  f$f�f(�fTPf/x�p  �8  f/hsgf/p��  f(�fY�f(�fY�f(- fY�fX-fY�fX- fY�fX-��Y�f(�f���X��Y��\Ń��f/`��   f(�fY�f(�fY�f(-�fY�fX-�fY�fX-�fY�fX-�fY�fX-�fY�fX-�fY�fX-�fY�fX-p�Y�f(�f���X��Y��\Ń���~�fW�f/XsO�~P�~-0�~��X�fs�,f��f~؍@�~,�h��~��\��Y��XH�^�f���   �~��~@�^�f��~�X��~$�`�f(�fY�f(�fY�f(- fY�fX-fY�fX- fY�fX-��Y�f(�f���X��Y��\��\��\�fVƃ��f/8u	f$���f/�sf$�Y҃��f$f`�Y҃���~��~@fT�f.�z�D$��f��X�`��ú�  ���T$�ԃ��T$�T$�$�~A  fD$���f�$�6F  �$�~$��ÍI �������̃��\$�D$%�  =�  u�<$f�$f��f���d$�n  f��f%�f-00f=��6  f��Y�f��-��X�f��\�f(��Y�fɁ�v ����?f(-������fY��\��Y��\�fxf����\�fY�f\�f(5��Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-��Y fX5�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��f��f%�f��f �\�f(�Ã�f�$�E  �$�~$����������̃��\$�D$%�  =�  ��  �<$f�$f��f����  f$f�f(�f(5�f(�f(�f��%�  ��@  +�-�<  Ё�   ��  fY�fX�f(�f\�fY�f(%�fY�f(-�f\�f~��ȃ�?������f\�f(��fY�f(�fY�fX��Y��X�f�fo5`f��fo5pf��fs�.fY��X�fV�f��X���~  ��|  w�Y��X�Ã���|$f�T$f�� f�$�,$����+�fo5Pf���  fn�fs�4fV���  fn�fs�4f$�$ft$�D$����f$$�$���$f$�l$��f�����  ���  s*�� t,��Á�   �r��+#��wr�$���9��s��ú   ��   ��fD$�T$�ԃ��T$���T$�$�|=  fD$�� �=  �s1�D$=   �sf �Y��   �f(�Y��   뙋$=  �w(�� u#�D$=  �uf���f��ú�  �]����D$%���=  �@�x���f$�X����f�$��C  �$�~$��Ã��\$�D$%�  =�  �8  �<$f�$f��f���#  f$fL$f=�Vf�VfT���fs�,f�� fV�f��%�   ��%�  �Y<�@f,�@�f(4�P"��  +у�ʁ�   ���  �    �� fn�f��fs����f(W��fs�&f�� fT%�V%�   ��%�  �Y�`*�Y,�`*�fX4�p.fV%�V�X�fT���fs�f�� f(W�\�f=0W%�  ��%�  �Y,��6�Y��6fX4Ő>fT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�f(Wf���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%(WfT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f(�N�Y��-��Y�f(�N�X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X�VfY��\�VfY��\�����f(��Nf(5 WfY�fX�fp���Y�fW���?  �X�f���X�f% Wfn��YT$�Y�fs�-fp�Df(=W�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��X��X��X��XÃ��fL$f�Vf~���fT�fs� f~Ɂ�  ���   ��� �B  �� �   �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$f(ѹ�  fn�fT�Vfs�4f��fPWf��fv�f��%�   �� ȁ�   ��r[�� f�Vf�V�5���f<$f(�f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=�Vf�V�Y�f~�fs� f~��� tRfT���fT�Vfs�,f�� fV�%�   ��%�  �Y<�@f,�@�f(4�P"�> �n����Ё������ u��T$��   ��� t0��#��  ��fn�fs� f�Vf$�^ʺ   �  ��#��� ��   fW����f�VfW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   umfL$f(ѹ�  fn�fT�Vfs�4f��f��f��fv�f��%�   =�   t-fL$f��% �  �� tfPW���fHW���fL$f��% �  �� �a  fW����fL$f��% �  �� �@  fW�����X��ĺ�  �  f$f~�fs� f~ҁ����¹    �� �k���f8WfpW�Yɺ   �Q  f$$fT$f�VfW�fT�fv�f��%�   =�   ��   f~��� u)fs� f~��  �?��   ��  �uf�V���f�VfW�fT�fv�f��%�   =�   ucf��f$$% �  ��  �у� ��   �� tf��%�  =�?  r!fW����f��%�  =�?  sfW����f@W����X��º�  �Vf~�fs� f~��������f�V�   �� t-f~�   %���=  �wr�� w���f@�   ��fD$�T$�ԃ��T$���T$���$�R4  fD$��(Ã� ~(=   �"  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X�V���� fY��\�VfY��\�����f(��Nf(5 WfY�fX�fp���Y��X��X�f% Wfnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(=W�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� A^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� � ������^�X��Y��Y��X�f��%�  �   =�  ������   �� ��������fhWfn��Y�fs�-fV��   �����   �� tfXW�Y`W�}���f`W�Y��l���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r�ɀ� fn�fs�-���f$$f�����  ���?  f��3�% �  �� �;����Y���f�$f�L$�9  �$�~$��Ã��\$�D$%�  =�  u�<$f�$f��f���d$�{  f��f%�f-00f=��6  f�_�Y�f�_�-��X�f�_�\�f(�_�Y�fɁ� v ����?f(-�_��W���fY��\��Y�_�\�fxf����\�fY�f\�f(5�_�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�_�Y fX5�_fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��,f��f=�u	�Y `�f�_�Y��\��Y�_Ã�f�$��9  �$�~$��ÍI �������̃��\$�D$%�  =�  ��   �<$�$������   f����%�  =�  t0��% �  u�Q����f�$�<$ uP�� �  uHf���� u>�ً���u$f��%��  uf��%��  uf�� %��  t�f�$�L$��  ��$    �D$  ���1   ���T$�ԃ��T$�T$�$�.  fD$���f�$�9  �$�~$��Ë��=�� �:  ���\$�D$%�  =�  u�<$f�$f��f���d$��9  � �~D$f(0`f(�f(�fs�4f~�fTP`f��f�ʩ   tL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$��-  ���D$��~D$f��f(�f��=�  |%=2  �fT `�X�f�L$�D$��``�f�@`fT `f�\$�D$���̃=�� ��9  ���\$�D$%�  =�  u�<$f�$f��f���d$��9  � �~D$f(�`f(�f(�fs�4f~�fT�`f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�,  ���D$��~D$f��f(�f��=�  |!=2  �fTp`�\�f�L$�D$����f��`fV�`fT�`f�\$�D$����������������WV�t$�L$�|$�����;�v;��h  �%L�s��  ���   ��  ��3Ʃ   u�%����  �%L� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����ȩ����   u������r*��$�ȩ��Ǻ   ��r����$�ܨ�$�ة��$�\����<�#ъ��F�G�F���G������r���$�ȩ�I #ъ��F���G������r���$�ȩ�#ъ���������r���$�ȩ�I ��������������|��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�ȩ��ة�� ��D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�d������$���I �Ǻ   ��r��+��$�h��$�d��x���Ī�F#шG��������r�����$�d��I �F#шG�F���G������r�����$�d���F#шG�F�G�F���G�������V�������$�d��I � �(�0�8�@�H�[��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�d���t�|������D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋T$�L$��t�D$�%L�s�L$W�|$��]�T$���   |�%����2  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�Q��`��3  Y�U��V��������EtV�+���Y��^]� U���   �} t��>  ��]ø����������Z������ �9��$��(����,�r��0����4����jh���pS  �E��uz�0G  ��u3��F  �B  ��u�,G  ����R  �������M  ���G  ��y��B  ���	J  ��x �/L  ��xj �iD  Y��u����   �I  �Ʌ�ue����~�H���e� �=�� u�D  ��B  �u��u�VI  �xB  �F  �E������   �   �u��u�=8��t�MB  ��p��u^�58���M  Y��u[h�  j�?Q  YY���������V�58���M  YY��tj V��@  YY����N��V�t  Y�������uj ��?  Y3�@�RR  � U��}u��K  �u�u�u�   ��]� jh����Q  3�@�u��u95���   �e� ��t��u5��`��t�uV�u�щE����   �uV�u�����E����   �]SV�u�������}��u(��u$SP�u����SW�u�������`��tSW�u�Ѕ�t��u*SV�u�������#��}�t��`��tSV�u�Ћ��}��E��������&�M�Q�0�u�u�u�   ��Ëe��E�����3��Q  �U��}u�uj �u�G����u�u�D=  YY]�U��} t-�uj �5������uV�n  ����P�s  Y�^]�U��V�u���woSW�����u�R  j��R  h�   �e@  ���YY��t���3�AQj P������u&j[9��tV�R  Y��u����  ���  ���_[�V��Q  Y��  �    3�^]����������̺����  ����<  �����������̃��\$�D$%�  =�  �  �<$f�$f��f����  f$f%pxf�xfW�fxx��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU�ofV�f($��`���X��\��Y��Y��Y����X��^�f=(xf-x�\�fs�?��fs�?�Y�fp�Df5 x�Y��Y�fW��Y��Y��X��Y��X�fp���X��X��Xă��-�  ��C�  �Y��\��Q�f��fs�fT=xfs���f%�x���\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<��o�Y�f(�w�Y��Y��\��X��\��X�f-x�\��X�f(x�^�f xf\��`���Y�%�   ���Y��Y��Y��Y��X�f���Y��X�f���X�fp���\��X�fVƃ���;  = 8  s]f�f(50xf�f(@xf(%PxfY�fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X����-�;  ���B  �Y��\��Q�f��fT= xfp�DfT x��f%�x���\��Y��X��Y��\����Y��Y��\��\��X��\�f(0xfp���\��X�fp���X��Y��X�fp���^�f(`xf(-@xf(PxfY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(�w�Y�fX�fp���Y�fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fVŃ���� = � ��   f~�fs� f~�����  �?+���� tpf$f~�fs� f~с��������  ��� }rfW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�@  fD$�� �fpxf�wf�w�X�fU�fV����f$fW��Xƺ�  �f$fW���f�����  �����  r�X�fV��Y����f�$�P  �$�~$��Ë������������̃��\$�D$%�  =�  �Y  �<$f�$f��f���D  f$�    f(�f�fs�4f�� f(�xf(yf(%�xf(5�xfT�fV�fX�f�� %�  f(��yf(��}fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(`yf(�f(pyfY�fY�fX�f(�y�Y�f(-�xfY�f(��xfT�fX�fX�fY��Y�fX�f(�f�fY�f(�fɃ��X��X��X��f$fW���� f�� �� wL���tb���  wpf$f(�xf(yfT�fV���� f�� �� t��fHyú�  �Ofy�^�f@y�   �4f0y�Y�������=��������  ���  s<fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$�b  fD$�� �f$f(�f~�fs� f~с��� ��� t���  �f�$��N  �$�~$�������Vjj �F  YY��V� ���������ujX^Ã& 3�^�jh���G  �e� �(:  �e� �u�#   Y���u��E������   ���G  Ëu��:  �U��QSV�5�W�5�����5���E��֋؋E�;���   ��+��O��rvP�O  ���GY;�sG�   ;�s�Ƌ]��;�rPS�sF  YY��u�F;�r>PS�_F  YY��t1��P��� �����u� ��K�Q� �����E�3�_^[��]�U���u�������Y���H]�U��U� ��ҋM#�#Mщ �]��O  ��tj�2O  Y� �t!j� �  ��tjY�)jh  @j�   ��j�'8  �U��E� �]�U���(  ��3ŉE��}�Wt	�u�R  Y������ ������jLj P�G�������������������0���������������������������������������������f������f������f������f������f������f��������������E�������E������ǅ0���  �@��������E�������E�������E������� ���������P��C  Y��u��u�}�t	�u�"Q  Y�M�3�_�������]�U��E�$�]�U���5$�����t]���u�u�u�u�u�   �3�PPPPP��������j�}�  ��tjY�)Vj� �Vj�s���V�NC  ��^�U��V�uWV�R  Y�N�����u�Y  � 	   �N ����  ��@t�=  � "   ��S3���t�^��t}�F�����N�F���^���F�  u*��P  �� ;�t�P  ��@;�uW�Q  Y��uV�\  Y�F  tz�V�+ʉM�B��FH�F��~QRW��Q  �����G�� �N�h���t���t�ǋ������������@��A tjSSW��Z  #����t%�N�E��3�@P�E�EPW�dQ  ����;]t	�N �����E��[_^]�U��V��M�F ��ufW�H1  ���~�Wl��Oh�N;��t�x��Gpu�^  ��F_;T�t�N�x��Apu�b  �F�N�Ap�u���Ap�F�
���A�F��^]� U���  ��3ŉE��E������SV�������EW�u�}������3��؉������������������������������������������������������������&  ����������������
  �@@ucP�O  Y�ȃ��t���t�������������@��B$��
  ���t���t�������������@��A$��T
  ���������F
  �3��������ȉ���������������������������������	  ������@����������	  �B�<Xw���������3����������ȁ�ǉ����������������������w	  �$�.�3���������؉������������������������������������<	  �� tF��t9��t/HHt���������	  ���������	  ����������  �����ˀ   ������*u/�������������������  ���؉������������  k�����
�����������  3��������  ��*u+������������������������p  ��������d  k�����
�����������>  ��ItE��ht8��������lt��w�,  ��   �����8lu@��   �������������� ������������ <6u�������4u�ǃ��� �  ����<3u�������2u�ǃ����������<d��  <i��  <o��  <u��  <x��  <X��  3��������3�������������P��P�hb  YY��t8������P�������������  ���������A���������������d  ������P�������������  ����  ��d��  �Q  ��S��   t|��AtHHtVHHtHH�  �� ǅ����   ��������������������@�   ���������������2  ǅ����   �  ��0  ��   ��   �������   ��0  u��   �������������������t�ʋ7����������  �S  ��u�5(�ǅ����   �ƅ�t3�If9t����u�+����<  ��X��  HHtp���'���HH�$  ����������  t0�G�Ph   ������P������P��b  ����tǅ����   ��G�������ǅ����   ��������  �����������t3�p��t,� ��   t�+�ǅ����   ���  3ɉ������}  �5$�V�`  Y�k  ��p��  ��  ��e�Y  ��g�K�����itd��nt%��o�=  ǅ����   ��y[��   �������M�����������`  ���  �������� tf���ǅ����   �z  ��@������ǅ����
   �� �  u��   ��  ���������3����  u��guVǅ����   �J;�~��������=�   ~7��]  W�;  ������������Y��t
���������
ǅ�����   ����������������������G�������������P��������������P������������VP�5(����Ћ�����   t!������ u������PV�54�����YY������gu��u������PV�50�����YY�>-�(�����   F����������ǅ����   j���s�����HH��������k  j'ǅ����   X���������|���Qƅ����0������ǅ����   �^�����3��������� t��@t�G���G����@t
�G���ȋ���O�����@t;�|;�s����߁�   �������� �  u����������y3�B�����   ������;�~�Ћ��u�������u��J�����������t=�������RPWQ�n_  ��0����������������9~������������N������밋������E�+�F��������   t6��t�>0t-N�������0�!��u�5$����I�8 t@��u�+Ɖ����������� ��  ��@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����������+���u������P������Wj �  ��������������������Q������P������P�  ����t��u������P������Wj0�  �������� ������t}��~y��H���������Pj�E􉍄���P������P��]  ����u?9�����t7������������P�������E�������P�t  ����������������u��(����������#������������Q������PV�:  ����������x#��t������P������Wj ��   ����������������tP����3�Y��������������������������������������������� _^[t
�������ap��M�3��6�����]��P  �    ���������_�g�����<�I�����U��U�B@t�z t/�Jx��M������ER��P�w���YY���u�E��]ËE� ]�U��V�u��~W�}W�uN�u�������?�t���_^]�U��V�uW�}��E�G@t� u
�M�E�N�& S�]��~@�EP�EKW� P�I����E���E�8�u�>*uPWj?�-����E����˃> u�E�[_^]��~$  ��u���Ã��U��V������MQ��    Y���   �0^]��J$  ��u���Ã��U��M3�;�0�t'@��-r�A��wjX]Í�D���jY;��#���]Ë�4�]�U��� �j�D��A  �u�v4  �=D� YYuj�A  Yh	 ��D4  Y]�U���$  j�A�  ��tjY�)�(��$�� ����5��=�f�@�f�4�f��f��f�%�f�-���8��E �,��E�0��E�<��������x�  �0��4��(�	 ��,�   �8�   jXk� ǀ<�   jXk� ���L�jX�� ���L�h$��������]�������U���0���S�ٽ\�����=|� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=|� t�#  ��8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����3  �   [�À�8�����=� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �H������������8�����s4�X��,ǅr���   �@������������0�����v�P�VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�X  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����K   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[��������̀zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����t����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-`���p��� ƅp���
��
�t���U��%H� ��S3�C	��j
���  ���L  3ɉH�3��V�5��W�}����_�O�W�E�M��E��ineI�E�5ntel�5��ȋE�5Genu���j�X��j Y���_�O�W�M�M�tC�E�%�?�=� t#=` t=p t=P t=` t=p u�=L����=L���=L��}�|5j3ɍu�X���Ƌ5���X�H�M��P�E�   t���=L��3���   tM���H�   �5����   t2��   t*���H�   �5��� t�� �H�   �5��_^3�[��]�U���(3��E��E�9P�t�5�����������E��   V;���  ��  ���  ��   jZ+���   H��   ����   H��   ����   HtN��	�#  �E�   �E���E�u� �E�]�� �E��]��P�]���Y����  ������ "   ��  �E���E�u�E�   � �E�]�� �E��]��P�]���Y�  �E�   �E����E����V  �U��E����l����E����;  �U��E����Q����E��놃�tfHtWHtHHt/���  ��	t���8  �E����   �E����   �E���E�u� ���   �E����   �E�   ������E�����   �E�   �E�������������   �$�s��E�����E�����E����E�$���E�,��u����E�4��i����E�<��]����E�D��E�u� �M��� �E�]�� �]��.�E�H����E�L����E�P��E�u� �E�]�� �]���E��E�   P�]���Y��u����� !   �E��^��]ð�����������d���B�6����$�-�����̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��R  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�R  ���$��X  �   ��ÍT$�mX  R��<$tmf�<$t�)X  =  �?s-����������������=� ��X  �   ����X  w8�D$��%�� D$u'��   ���t���������W  ���� u�|$ u����-`��   �=� �*X  �   ����3W  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��X  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�X  ���$�rW  �   ��ÍT$�W  R��<$t6f�<$t�-x�����=� �PW  �   ����MW  ��V  �&��� u�|$ u����-j��   �t���뻸   �=� �W  �   ����V  Z������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�Z  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�UZ  ���$�RV  �   ��ÍT$��U  R��<$tPf�<$t�-x�������z�=� �,V  �   �С�)V  �-z���������z��������U  ���� u�|$ u����-`��   �=� ��U  �   �С��T  Z�������̃=�� tn���\$�D$%�  =�  u�<$f�$f��f���d$uA�-[  ��=�� t<���\$�D$%�  =�  u�<$f�$f��f���d$u��Z  ����9�������c�������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uZ�Z_  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�_  �����$�T$�D$�   ��ÍT$�8T  ��P��<$f�<$t��S  ��  ��T$��  ���   �	T  ��   �  ���   �L$���S  ���S  ��u���=� �)T  ���   �dT  �=� �T  ���   ��R  ZÍT$�S  �D$uA�3���   ���D$u����   �3��3�%�� D$uÍT$�[S  �D$��%  ����� =  �uT$u���u���t��Q���$�\$��q�i  ��Y�a���t���eS  �   �B����D$%�� D$������؋D$%���D$t=�f   �l$���D$�   t�-����t��   ���������S  ����R  ������R  ���   ��������������-`��   ���������ٱ ����u���������ٛ���u�����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��i  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�ui  ���$�R  �   ��ÍT$�Q  R��<$tPf�<$t�-x�������z�=� ��Q  �   ����Q  �-z���������z��������?Q  ���� u�|$ u����-`��   �=� ��Q  �   ���P  Z�������̃��$�MQ  �   ��ÍT$��P  R��<$�D$tQf�<$t�P  �   �u���=� �#Q  �   � �� Q  �  �u,��� u%�|$ u���P  �"��� u�|$ u�%   �t����-`��   �=� ��P  �   � ���O  Z�j
���  ���3��U��QQSV���  V�5��r  �E��YY�M��  ��#�QQ�$f;�uT�q  YY��~-��~��u#�ESQQ�$j�Pl  ���qVS�Jr  �EYY�c�E���S�����\$�$jj�?�0i  �U��E��������DzV��S���r  �E�YY��� u�S�����\$�$jj�7i  ��^[��]�U��QQSV���  V�5���q  �E��YY�M��  ��#�QQ�$f;�uT�p  YY��~-��~��u#�ESQQ�$j�yk  ���qVS�sq  �EYY�c�E���S�����\$�$jj�?�Yh  �U��E��������DzV��S���.q  �E�YY��� u�S�����\$�$jj�`h  ��^[��]Å�uf���fn�f`�fa�fp� SQ�ك���ux�ڃ���t0ffAfA fA0fA@fAPfA`fAp���   KuЅ�t7����t��I f�IKu���t����t
f~�IJu���t�AKu�X[��ۃ�+�R�Ӄ�t�AJu���t
f~�IKu�Z�^���̋T$�L$��   u@�:u2��t&:au)��t��:Au��t:au������uҋ�3���������Ë���   t���:u����t���   t�f���:u΄�t�:auń�t����jh���   j�p  Y�e� �u�F��t0�X��T��M��t9u,�A�BQ�,���Y�v�#���Y�f �E������
   �   Ë���j�q  Y�U��j �u�u�u�u�u�u�   ��]�U��E��et_��EtZ��fu�u �u�u�u�u��  ��]Ã�at��At�u �u�u�u�u�u�}  �0�u �u�u�u�u�u�   ��u �u�u�u�u�u��  ��]�U���,SVWj0X�u���E��  �M�3ۍM������}��y���u��t�M��u	����j��G�;�w����j"_�8�������  �U��Z�E����%�  =�  uy3�;�uu���;�t�A�j WP�^SR��  ������t� �  �;-u�-F�}��j0X�����$�x�F�FjeP��y  YY��t�����ɀ����p��@ 3��O  3���   ��t�-F�} �]j0X�����$�x�ۈF�Jۃ����  ���'3���]�u'j0X�F���B�
%�� �u3��E���E��  ��F1����F�M��u� ��Eԋ��   � � ��B%�� �E�w	�: ��   �e �   �E��M��~S��R#E#ыM����� ���A~  j0Yf�����9vËM�U�F�E���E�E�����O�M�E�f��y�f��xW��R#E#ыM����� ����}  f��v6j0�F�[���ft��Fu�H��]�;E�t���9u��:��	�����@���~Wj0XPV���������E�8 u���} �4�U����$�p���R�q}  �ȋ�3����  #�+M��x;�r	�F+����F-��������0��;�|A��  ;�rPRSQ�C|  0�U�F3�;�u;�|��drPjdSQ� |  0�U�F3�;�u;�|��
rPj
SQ��{  0�U�F�]�3���0����F�}� t�M܃ap���_^[��]�U��j �u�u�u�u�u�V  ��]�U����M�SW�u �5����]��t�} w	�K���j��U3����ǃ�	9Ew�-���j"_�8�q�����   �} t �M3�����P3��9-���P��  �UYY�EV��8-u�-�s��~�F�F�E����   � � �3�8E�������9Et��+�Ehh�PV��j  ����uv�N9}t�E�U�B�80t-�RJy���F-jd[;�|��� Fj
[;�|��� F V���^t�90uj�APQ�o  ���}� t�M��ap���_[��]�WWWWW�~����U���,��3ŉE��E�M�S�]VW�}j^VQ�M�Q�p�0�y  ����u������0�(������t�u��u
�����j^����;�t3��΃}�-��+�3�����+ȍE�P�CPQ3Ƀ}�-��3�������P�nv  ����t� ��u�E�j P�uSVW��������M�_^3�[�2�����]�U����E�M�SV�u�@H�E������u��t�} w�"���j[��f����   3�W�}8]t�M�;�u�U3��:-���f�00 �E�8-u�-F�@��jV�  Y�0FY����~JjV�  �E�YY���   � � �F�E�@��y&8]t�������;�|��WV�l  Wj0V�������_�}� t�M�ap�^��[��]�U���,��3ŉE��E�M�SW�}j[SQ�M�Q�p�0��w  ����u�+�����r������lV�u��u������Z������S���;�t3��΃}�-��+ȋ]�E�P�E��P3��}�-Q���P�t  ����t� ��u�E�j PSVW�g�����^�M�_3�[腞����]�U���0��3ŉE��E�M�SW�}j[SQ�M�Q�p�0�!w  ����u�j�����������   V�u��u�O�����������   �E�3�H�}�-�E�������9;�t��+��M�Q�uPS��s  ����t� �S�E�H9E������|+;E}&��t
�C��u��C��u�E�jP�uVW��������u�E�jP�u�uVW�I�����^�M�_3�[膝����]�U��j �u�   YY]�U���W�u�M��Z����U�}��
��t���   � � :�tB�
��u��B��t4�	<et<EtB���u�V��J�:0t����   ��:uJ�BF���u�^�}� _t�E��`p���]�U��j �u�u�u�   ��]�U��QQ�} �u�ut�E�P�t  �M�E���E��A��EP�t  �M�E�����]�U��j �u�   YY]�U����M�V�u�o����u�P�j  ��e�F�P�Bi  ��Yu��P�j  Y��xu���E�����   � � �F���ȊF��u�^8E�t�E��`p���]�U��E�������Az3�@]�3�]�U��W�}��tV�uV��8  @P�>VP�\j  ��^_]�Vh   h   3�V�!v  ����u^�VVVVV�+����V3����� ��������(r�^�U��V��  �����E  �V\��W�}99t�����   ;�r�   ;�s99t3Ʌ��  �Q���  ��u�a 3�@��   ��u�����   �ES�^`�F`�y��   j$_�F\�d �����   |�9�  ��~du�Fd�   �   �9�  �u	�Fd�   �u�9�  �u	�Fd�   �d�9�  �u	�Fd�   �S�9�  �u	�Fd�   �B�9�  �u	�Fd�   �1�9�  �u	�Fd�   � �9� �u	�Fd�   ��9� �u�Fd�   �vdj��Y�~d�	�q�a ��Y�^`���[�3�_^]�U��csm�9Eu�uP����YY]�3�]�jh ��J  �u����   �~$ t	�v$�}���Y�~, t	�v,�n���Y�~4 t	�v4�_���Y�~< t	�v<�P���Y�~@ t	�v@�A���Y�~D t	�vD�2���Y�~H t	�vH�#���Y�~\p�t	�v\����Yj�/c  Y�e� �Nh��t�����u��0�tQ�����Y�E������W   j��b  Y�E�   �~l��t#W�e-  Y;=��t����t�? uW��+  Y�E������   V����Y�  � �uj�d  YËuj��c  Y�U��8����t'V�u��uP�l  ��8�Yj P�{  YYV����^]�V�   ����uj�  Y��^�VW���58����$  ��Y��uGh�  j�  ��YY��t3V�58��  YY��tj V�%   YY���N���	V����Y3�W�$�_��^�jh(��X  �u�F\p��f 3�G�~�~pjCXf���   f���  �Fh0����   j�a  Y�e� �Fh�����E������>   j�la  Y�}��E�Fl��u����Fl�vl��)  Y�E������   �  �3�G�uj�b  Y�j�b  Y��  �Jb  ��u�c   3��h:��  �8�Y���t�Vh�  j�T  ��YY��t-V�58���  YY��tj V�����YY���N��3�@^��   3�^á8����tP�r  �8��Y��`  U��Q�E�Ph�j �,���th(��u��0���t�u�Ћ�]�U���u�����Y�u�(��VW�5�����5p�����t�> t�6�����Y��u�5p�SV�����5l�3ۉp�Y��t9t�6�ɾ��Y��u�5l�V跾���5h��l�覾���5d�蛾������h����d�;�t9��tW�w���YV� ���������tP�[���Y��������tP�E���Y����T���0N[u�T��0�;�tP����Y�5T�_^�U����  �u�;  Yh�   �   �jj j �>  ���U��=�` th�`�fp  Y��t
�u��`Y����h�h���   YY��uChd�����$ �h���v   �=�� YYth���p  Y��tj jj ���3�]�U��j j�u�   ��]�Vj � ���V�  V�����V����V�  V��p  V��p  ��^��	  U��ESV�u3�+ƃ���9uW���#�v���t�Ѓ�C;�r�_^[]�U��V�u3����u���t�у�;ur�^]�j��]  Y�j�@_  Y�jhP��V  j��]  Y�e� �=\���   ���   �E����} ��   �5���5��֋؉]ԅ�tt�5���֋��]�}��}܃��}�;�rWj � �9t�;�rG�7�֋�j � �����5���5��։E��5���֋M�9M�u9E�t��M�ى]ԉE����h0�h �����YYh8�h4�����YY�E������    �} u)�\�   j�-^  Y�u�^����} tj�^  Y��y  ��<�3ɣ��������Ã%�� �jdhp��
  j�u\  Y3ۉ]�j@j _W��
  YY�ȉM܅�uj��E�Ph���]  ������[  ����=��   ;�s1f�A 
�	��Y�a$��A$$�A$f�A%

�Y8�Y4��@�Mܡ���ƍE�P�L�f�}� �/  �E����$  ��M���E���E�   ;�|�ȉM�3�F�u�9��} j@W�
  YY�ȉM܅���   ����M���}�j�[�E؋U�;���   �2���t[;�tW� �tQ�uV�D��U���t<����������4����u܋��E؊ �Fj h�  �FP�V  ���F�U��M�G�}ԋE�@�E؃��U�냉���=������   ;�s$f�A 
�	��Y�a$�f�A%

�Y8�Y4��@�M���F�uЋM�� ���j�[3��}ԃ���   ����5���u܃>�t9t�F��F�   �F���uj�X�
�G�������P�@��E���tL��tHP�D���t=�M�%�   ��u�F@���u	�F�Fj h�  �FP�J  ���F��F@�F������t���XG�=����]��   3��	  �j�@[  Y�VW����>��t7��   ;�s"���� tW�H����@��   �G�;�r��6�n����& Y������|�_^�U��QQ�=�� u�\%  SVWh  ���3�WS����P��5���=t���t8u���E�P�E�PSSV�]   �]��������?sE�M����s=��;�r6R�  ��Y��t)�E�P�E�P��PWV�    �E���H�=d��`�3�����_^[��]�U��ES�]V�uW�# �}�    �E��t�8���E3ɉM�>"u3�����F�Ȱ"�M�5���t��G�F�E��P�{k  Y��t���t��GF�E��t�M��u�< t<	u���t�G� �N�e �> ��   �< t<	uF��> ��   �U��t�:���U�E� 3�B3��FA�>\t��>"u3��u�} t�F�8"u���3�3�9E���E���I��t�\G���u���tA9Mu< t8<	t4��t*��P�j  Y��t��t��GF���G���tF��F�o�����t� G��-����U_^[��t�" �E� ]Ã=�� u�2#  V�5�W3���u����   <=tGV�R*  FY����u�GjP�x  ���=l�YY��tʋ5�S�> t>V�*  �>=Y�Xt"jS�G  �YY��t@VSP�yV  ����uH���> uȋ5�V苵���%� �' 3����   Y[_^��5l��e����%l� �����3�PPPPP�=����U����e� �e� ��VW�N�@��  ��;�t��t	�У��f�E�P�\��E�3E�E���1E��X�1E��E�P�T��M��E�3M�3M�3�;�u�O�@����u��G  ��ȉ��щ�_^��]�U��QW�`���3���tuV��f9t��f9u���f9u�SPPP+�P��FVWPP�8��E���t7P�;  ��Y��t*3�PP�u�SVWPP�8���u	S�A���Y3�W�d����	W�d�3�[^_��]�U�� �3�t�u��]�]�%��U���3��ut��]����]�U���3��ut��]����]�U���3��u�ut��]����]�U���3�t�u�u�u��]��u�u�p�3�@]�U��QV�5����y%�t�3�3��u�tV�M�Q�Ѓ�zuF�5��3���^����]���VWh8�����50���hT�W��3�h`�W� ���3�hh�W����3�ht�W����3�h��W����3�h��W����3�h��W����3�h��W����3�h؜W����3�h�W� ���3�h�W�$���3�h$�W�(���3�h<�W�,���3�hT�W�0���3�hh�W�4���3��8�h|�W��3�h��W�<���3�h��W�@���3�hԝW�D���3�h��W�H���3�h�W�L���3�h$�W�P���3�h8�W�X���3�hH�W�T���3�hX�W�\���3�hh�W�`���3�hx�W�d���3�h��W�h���3�h��W�l���3�h��W�p���3�h̞W�t���3��x�hܞW��3�h��W�|���3�_���^�U���u�t�]�U���u�x�P�|�]�U��j �l��u�h�]�U��VW3�j �u�u�Oe  ������u%9��vV�������  Y;5��v������uŋ�_^]�U��SVW�=��3��u�K�����Y��u#��tV�X����=�����  Y;�v������u�_^��[]�U��VW3��u�u�d  ��YY��u*9Et%9��vV�������  Y;5��v������uË�_^]�VW�p��p�����t�Ѓ�;�r�_^�VW�x��x�����t�Ѓ�;�r�_^�������������h�d�5    �D$�l$�l$+�SVW��1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q��������U���S�]VW�E� �{�s3=��E�   ����t�O�30�$����G�O�30�����E�@f��   �E�E�E�E�C��C�E������   �@�@�L�����E���t{���R  ��M����~   ~h�E�8csm�u(�=�� th����`  ����tj�u������U�M��Q  �E�U�9Pth�V����Q  �E�X����tu�f�M��]��Ã���^�����tG�!�E�    ��{�t6h�V�˺�����Q  ����t�O�30�����W�O�32������E�_^[��]ËO�30�����G�O�30�Մ���M��֋I�Q  �U���5������t�u��Y��t3�@]�3�]�U��E���]�j�)d  Y��tj�d  Y��u�=��uh�   �1   h�   �'   YY�U��M3�;��t
@��r�3�]Ë��]�U����  ��3ŉE�V�uWV������Y���y  Sj�c  Y���  j�c  Y��u�=����   ���   �A  h��h  h���,b  ��3ۅ��1  h  h��Sf��������  ��uh�Vh����a  ������   h���6b  @Y��<v5h���%b  jh��El���-����+�VQ�b  ������   h$�h  ���V�a  ������   Wh  V�a  ����u}h  h0�V��b  ���Wj��@�����tI���tD3ۋˊO�����f9Ot	A���  r�S������]�P�����P�  YP�����PV���[�M�_3�^艂����]�SSSSS����������������������7   ���"�.   ��������2��ƅp��������������
�t����
�t�����������������������ݽ`������a���u2����X��������-j����
�t����
�t�������
�t�����������؊�� ����������������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�Yc  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�c  ���$��'  �   ��ÍT$�'  R��<$tmf�<$t�I'  =  �?s+��������������=� ��'  �   ����'  w:�D$��%�� D$u)��   ����-j�t�����'  ���� u�|$ u����-`��   �=� �J'  �   ����S&  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�g  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�Eg  ���$�&  �   ��ÍT$�=&  R��<$tL�D$f�<$t�-x��  �t^�   �uA������=� �\&  ����   �Y&  �   �u�ԩ�� u�|$ u%   �t����-`��   �"�%  ���� uŃ|$ u����-���   �=� ��%  ����   ��$  Z�U���uj �u�u�u�   ��]�U��� �e� 3�W�}�jY�9Eu�����    �G�������x�EV�u��t��u������    �#�������S�����M�;�w�E��u�E��E�B   �u�u��u�u�P����������t�M�x�E��  ��E�Pj �
���YY��^_��]�U��} u�i����    謲�����]��uj �5�����]��5�����U��E������������]�j$h���3����e� �e� 3ۉ]�3��}؋u��Pt��jY+�t"+�t+�t^+�uH�*������}؅�u����b  �E�������^�w\V�Q  YY���E� �V�ƃ�t6��t#Ht�����    �ֱ����E��������E��������E������3�C�]�P���E܃���   ��uj�D�����tj ��F  Y�e� ��t
��t��u�G`�Eԃg` ��u?�Gd�E��Gd�   ��u-���щU̡��;�}$k��G\�d B�Ű���j � ��M��E������   ��u �wdV�U�Y��u�]��}؅�tj �G  Y�V�U�Y��t
��t��u�EԉG`��u�EЉGd3�������U��U� �V�u9rtk���E;�r�k�M;�s	9ru���3�^]�U��E��t���8��  uP�{���Y]�U��SVW3���   �;�+���jU�4���u�   ����ty�^���~;�~Ѓ�������_^[]�U��} t�u����Y��x=�   s	��Щ]�3�]�U��p�3�t3�QQQ�u�u�u�u�u�u��]��u�u�u�u�u�u����YP���]�U��V�u3���t^�MSW�}jA[jZZ+��U�jZZ�f;�rf;�w�� ������f;�rf;Ew�� ����Nt
f��tf;�t�����_+�[^]Ã%�� á��Vj^��u�   �;�}�ƣ��jP�������YY��ujV�5���������YY��ujX^�3ҹ����� �R��(�}�����3�^��me  �=�� t�d  �5��譢���%�� Yø���U��V�u���;�r"���w��+�����P�C  �N �  Y�
�F P���^]�U��E��}��P�qC  �EY�H �  ]ËE�� P���]�U��E���;�r=�w�`���+�����P�D  Y]Ã� P���]�U��M�E��}�`����AP�gD  Y]Ã� P���]�U��E��u�K����    莭�����]Ë@]�U��M���u�&���� 	   �8��x$;��s�������������D��@]������ 	   �4���3�]�jh�������3ۉ]�u���u萻���轻��� 	   �   ����   ;5����   ���������������D8��u
�G����  �jV�rd  Y�e� �����D8t�u�uV�^   ������E���� 	   �����  ����}��E������
   ���(�u�}�V�e  Y��ں�������� 	   �J�������[����U���  ��f  ��3ŉE���D��� �E�MV3���8���W3���0�����@���9uu3��  ��u�n���!0蛺���    �ޫ�������  �Ћ���������(���S������$����\$�����t��u+�E�Шu����!0�@����    胫���  ��8����D tjj j P�  ����8��������Y���P  ��(�����$��������D��2  ����3ɋ@l9��   �����P��(�������<�����$��������4�������  9�<���t����  �����0���3�!�8����������4�����,���9M��  ��,���3҉�@���ǅ���
   !�<�������  �3���$�����
���������(���������<���9|8t�D4�E�<����U�j!|8�E�P�Z��P�  Y��tD��0�����,���+�E����  jR��4���P�Od  ������  ��,���@��@����&j��,�����4���P� d  �������  ��,���3�@��@���QQj��,����E�Pj��4���PQ������8���<�������  j ��8���Q��$���P�E�P��(��������4������L  ��@�����D����<���9�8����I  9����tK��$�����8���j Pj�E��E�P��(��������4�������   ��8�����  ��D���F��4����   ��t��u3�3�f;������4�������<�����@�������,�����@�����t��uKQ��b  Y��4���f;�uu��9�<���t"jXP��4�����b  Y��4���f;�uOF��D�����@�����,���;U������E  ��(���F���$��������D
4�����D8   �  �����
  ��(���������$����D��u  ��0���3���4������  �]��8�������  3ɍ�������<���+�0���;�sD�
B@�������
��8�����<���u��D����GA������G��8���A��<������  r���$���������+��� ���j PW������P��(��������4���������� ���9� ���|��8�����+�0���;��A�����4�����D�������  ����  j[;���  耵��� 	   �A������  �ʀ���   9u�|  ǅ���
   ����� ��������j+����^;Es3�9����f;����u��D���f�3����f�;�������  rȍ�������<�����$���+�j �� ���PS������P��(��������4�����@�����4����������� �����@���9� ����������<�������0���+�;E�.���������]��8�������  ǅ���
   ����� ��H�����8���+ʋ����;�s;�7������8���f;����uj_f�8����8�����f�0�������  r�3�������VVhU  Q��H���+��+���P��PVh��  �8���@�����4�����<������ ���3ɉ�@���j +��� ���RP���������$���P��(��������4�����t��@���� �����<�����@���;�������@�������<�����4���;��������8�����0���+�@���;�������w���j �� ���R�u��0����4������=����� ���3��G���W�Ʋ��Y�<��0�����(�����$��������D@t	�:u3��趲���    �w����  ����+��[�M�_3�^�oo����]�jhЗ��������u؉u܋}���u�8����  �d���� 	   �   ����   ;=����   �����E�߃��������D��tpW� [  Y�e� �E�����Dt�u�u�uW�g   ������������ 	   謱���  �މu؉]��E������   ���+�}�]܋u�W�3\  Y��{����  觱��� 	   �����֋�������U��QQV�uWV�[  ���Y;�u�u���� 	   �ǋ��D�u�M�Q�u�uP�����u��P�$���Y�Ӌƃ����������d0��E��U�_^��]�U�����V�   V�O���Y�M�A��t	�I�q��I�A�A�A   �A�a �^]�U��U3�SVAW�����rx��t�������   ��t�����r|��t�������   ��t����j�r[�~�T�t�>��t�����~� t�~���t������Kuҋ��   �   ��A_^[]�U��SV�u3�W���   ��tf=خt_�Fx��tX9uT���   ��t9uP�w������   �+\  YY�F|��t9uP�Y������   �	]  YY�vx�D������   �9���YY���   ��tD9u@���   -�   P�������   ��   +�P�������   +�P��������   ���������   =X�t9��   uP��\  ���   �Ô��YYjX���   �E�~��T�t���t�8 uP蘔���3葔��YY�E�� t�G���t�8 uP�t���Y�E����H�Eu�V�^���Y_^[]�U��U����   SV���W�����Jx��t�������   ��t�����J|��t�������   ��t����j�J[�y�T�t�9��t�����y� t�y���t������Kuҋ��   ���   ��1N_^[��]�jh��`����e� �l������x��Npt"�~l t�T����pl��uj �j���Y���n����j�4  Y�e� �5���FlP�!   YY���u��E������   뼋u�j��5  Y�U��W�}��t;�E��t4V�0;�t(W�8�����Y��tV�����> Yu����tV�F���Y��^�3�_]Ã=�� uj��M  Y���   3��U��E-�  t&��t��tHt3�]á��]á��]á��]á��]�U����M�j �����%� �E���u��   ����,���u��   �������u�E���   �@�}� t�M��ap���]�U��S�]VWh  3��sWV�����{3��{����  �  �{����0�+��7�FIu���  �   �9�AJu�_^[]�U���   ��3ŉE�SV�u������WP�v�İ3ۿ   ����   �È�����@;�r�����������ƅ���� ��Q���;�sƄ���� @;�v�����u�S�v������PW������PjS�`  S�v������WPW������PW��  S�^  ��@������S�vWPW������Ph   ��  S�^  ��$����M�����t�L��������t�L ��������  ���  A;�r��Yj���  ��X+������������� ��w
�L�A �������w��H �A������������  A;�r��M�_^3�[�g����]�jh������3��u���������x��Opt9wlt�wh��uj �����Y��������j�1  Y�u��wh�u�;5T�t4��t�����u��0�tV�Ï��Y�T��Gh�5T��u�3�@���E������   둋u�j�"2  Y�jh0��8�������E����؉]��<����sh�u�����Y�E;F�h  h   �'���Y�؅��U  ��   �E��ph���3��3S�u�A  YY���}���  �E��Hh�����u�Hh��0�t
Q�����Y�E��Xh3�@���E��@p��   �x���   j��/  Y�u��C����C�����  ���ΉM��}f�DKf�M �A��ΉM��  }�D��(�A��u��   }��  ��0�F��T������u�T�=0�tP�=���Y�T�3�@���E������   �1�}j�0  Y��#���u��0�tS� ���Y茨���    �3���������U��� ��3ŉE�SV�u�u�6�����Y��uV����Y3��  W3��ϋǉM�9�X���   A��0�M�=�   r����  ��   ����  ��   ��P�������   �E�PS�İ����   h  �FWP�J����^��3ۉ�  C9]�vO�}� �E�t!�H��t�����LA;�v����8 uߍF��   �@Iu��v�"�������  �^��~3��~����   9=�tV�����   ����   h  �FWP譈����kE�0�E���h��E�8 ��t5�A��t+������   s��P�DB�A;�v���9 u΋E�G���E��r�S�^�F   �o�������  �E��Nj��\�_f��Rf��IOu�V�I���Y3�_�M�^3�[�pc����]�U����u�M��V����E�ȋE����   �H% �  �}� t�M��ap���]�U��j �u����YY]������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�3���9����U���S�]W�}��u��t�E��t�  3���E��t��V�����v�b���j^�0視���X�u�M��#����E�3�9��   ubf�E��   f;�v;��t��tWVS蒆��������� *   �����0�}� t�M��ap���^_[��]Å�t��t_��E��t��    �эM�uQVWSj�MQV�p�8��ȅ�t9uu��E��t�������zu���t��tWVS������艤��j"^�0�͕���o���U��j �u�u�u�u�������]��V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� S��QQ�����U�k�l$���   ��3ŉE��CV�sW���|����Ht+Ht$HtHtHtHHtHuzj��   �nj�
j�j�j_Q�FPW�!  ����uG�K��t��t��t�e����E��F�����]��E��FP�FPQW��|���P�E�P� #  ����|���h��  Q�(  �>YYt�=|� uV����Y��u�6��%  Y�M�_3�^�_����]��[���U�������$�~$�   ��fD$f% �f0�fW�f(���fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU`�fV�f($�`����X��\��Y��Y��Y����X��^�f��f-���\�fs�?��fs�?�Y�fp�Df5���Y��Y���fW��Y�f\%`��Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<�`��Y��Y��Y��\�fTp��X��\��X�f-���\��X�f���^�f��fX�`����Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(5��f�f(��f(% �fY�f(-`���fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT= �f%8�f(���Y�f(���\�f( �fp�D�Q�fY�fp�Df��fY�fX�f��fY�����Y�fX�fp�D�Y�fTp�fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�P���fD$����fD$�D$���f������fn�fp� f��f��fT�fT��X�fD$�D$���f`�fh��X�fD$�D$���fW��Xƺ�  �J���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�U������E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��p��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z����������������������   s��������������������������   v���������U�������$�~<$�   ���~|$f�f(�fT��f/����  �U  f/��snf/����  f(�fY�f(�fY�f(-��fY�fX-��fY�fX-��fY�fX-p��Y�f(�f���X��Y��\�f�|$�D$�f/����   f(�fY�f(�fY�f(-`�fY�fX-P�fY�fX-@�fY�fX-0�fY�fX- �fY�fX-�fY�fX- �fY�fX-���Y�f(�f���X��Y��\�f�|$�D$��~�fW�f/��sO�~���~-���~��X�fs�,f��f~؍@�~,�h��~��\��Y��X���^�f���   �~��~���^�f��~�X��~$�`�f(�fY�f(�fY�f(-��fY�fX-��fY�fX-��fY�fX-p��Y�f(�f���X��Y��\��\��\�fV�f�D$�D$�f/��u�D$�f/ �s�������$�$���D$������D$��~��~��fT�f.�z�D$��������ú�  ���T$�ԃ��T$�T$�$��������D$Ð����U�������$�~$�   ��fD$f��f%�f-00f=��B  fP��Y�fX��-��X�fp��\�f(`��Y�fɁ�v ����?f(-@������fY��\��Yx��\�fxf����\�fY�f\�f(5 ��Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-0��Y fX5�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f���\�fL$�D$��������I ����U�������$�~$�   ��fD$f�f( �f(5 �f(0�f(@�f��%�  ��@  +�-�<  Ё�   ��(  fY�fX�f(�f\�fY�f(%P�fY�f(-`�f\�f~��ȃ�?������f\�f(�p�fY�f(�fY�fX��Y��X�f�fo5��f��fo5��f��fs�.fY��X�fV�f��X���~  ��|  w�Y��X�fD$�D$��Ã���|$f�T$f�� f�$�,$����+�fo5��f���  fn�fs�4fV���  fn�fs�4f$�$ft$�D$����f$$�$���$f$�l$��f�����  ���  s'�� t)�Z��   �r��+#��rJw�T$���9��r<��   ��   ��fD$�T$�ԃ��T$���T$�$����fD$����fD$�D$���=  �s1�D$=   �sf���Y��   �f���Y��   뉋T$=  �w�� u�D$=  �u�������ú�  �V����D$%���=  �@s�fD$�Xp���fD$�D$��ÍI ƅp����
�u;�����ƅp����2������+  ������a���t������@u��
�t���Ҙ���F  �t2��t��������Ș���^��������-��ƅp����������ݽ`������a���Au����ƅp������-���
�uS��������
�u�����n�����   ����
�u���u
�t���ƅp����-����u�
�t��������-������Ș��X��ݽ`������a���u���-��
�t���ƅp�������������-��ƅp����
�u����-��������-���ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u����������ٛ���t�   ø    ���   ��V��t��V���$���$��v��  ���f���t^��t��������������U���������$�\$�   ��fD$f=�.f�.fT���fs�,f�� fV�f��%�   ��%�  �Y<� �f,� ��f(4�0���  +у�ʁ�   ���  �    �� fn�f��fs����f/��fs�&f�� fT%�.%�   ��%�  �Y�@�Y,�@�fX4�PfV%�.�X�fT���fs�f�� f/�\�f=/%�  ��%�  �Y,�`�Y�`fX4�pfT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�f/f���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%/fT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f(�&�Y��-��Y�f(�&�X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X�.fY��\�.fY��\�����f(��&f(5�.fY�fX�fp���Y�fW���?  �X�f���X�f% /fn��YT$�Y�fs�-fp�Df(=�.�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��XŃ��X��X��X�fD$�D$���fL$f�.f~���fT�fs� f~Ɂ�  ���   ��� �  �� �  �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$fT$��  fn�fT�.fs�4f��f0/f��fv�f��%�   �� ȁ�   ��r^�� f�.f�.�&���f|$fd$f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=�.f�.�Y�f~�fs� f~��� tRfT���fT�.fs�,f�� fV�%�   ��%�  �Y<� �f,� ��f(4�0��> �\����Ё������ u��T$��   ��� t1��#��  ��fn�fs� f�.fT$�^ʺ   �  ��#��� ��   ���f�.fW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   uefL$fT$��  fn�fT�.fs�4f��f��f��fv�f��%�   =�   t#fL$f��% �  �� t�0/��(/�fL$f��% �  �� �G  ���fL$f��% �  �� �+  ����X��ĺ�  �  fT$f~�fs� f~ҁ����¹    �� �����f/fP/�Yɺ   �H  fd$fT$f�.fW�fT�fv�f��%�   =�   ��   f~��� u fs� f~��  �?��   ��  �u���f�.fW�fT�fv�f��%�   =�   uUf��fd$% �  ��  �у� ��   �� tf��%�  =�?  r���f��%�  =�?  s���� /��X��º�  �cf~�fs� f~��������f�.�   �� t:f~�   %���=  �w%r�� w��fD$�D$���f ��   ��fD$�T$�ԃ��T$���T$���$�����D$��Ã� ~(=   �<  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X�.���� fY��\�.fY��\�����f(��&f(5�.fY�fX�fp���Y��X��X�f% /fnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(=�.�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� N^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� ������fD$�D$���^�X��Y��Y��X�f��%�  �   =�  ������   �� �������fD$�D$���fH/fn��Y�fs�-fV��   �����   �� tf8/�Y@/�e���f@/�Y��T���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r �ɀ� fn�fs�-��fD$�D$���fd$f�����  ���?  f��3�% �  �� �-����K�����$    ��$    �U��QQ�EQQ�$�.;  YY��uJ�EQQ�$�C  �E����YY����Dz+���QQ�U��$�   �E�����YY��DzjX�	3�@���3���]�U���E�  �V3���  ��9Mu:9uu|��������z�����h���   ��������A�E��   ������   9EuB9uu=��������z�������   ������A�Eu�h��   �p�3��F�   ��9Mu-9u��   ���E������A�m����������E{[�����U9Eu]9uuX�EQQ�$�������EYY�ы�����Au�����h���u���������z��u������E��	�M�������^]���U�������$�~$�   ��fD$f��f%�f-00f=��B  f�7�Y�f�7�-��X�f�7�\�f(�7�Y�fɁ� v ����?f(-�7�`/���fY��\��Y�7�\�fxf����\�fY�f\�f(5p7�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�7�Y fX5`7fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y�7fD$�D$���f�7�Y��\��Y�7fD$�D$����ؔ���U��QQ�E���]��E���]�U��E� tj��t3�@]ètj��tjX]������]�S��QQ�����U�k�l$���   ��3ŉE�V�s �CVP�s�   ����u&�e��P�CP�CP�s�C �sP�E�P�  �s ���s�c����=|� Yu)��t%�CV���\$���\$�C�$�sP�  ��$�P�X  �$��  V��  �CYY�M�3�^�?����]��[�U���S�]V�����t�Etj��  Y����  ��t�Etj��  Y����u  ����   �E��   j�  �EY�   #�tT=   t7=   t;�ub�M������x���{L�H�M�������{,�x��2�M�������z�x���M�������z�h���h���������   ����   �E��   W3���tG�M���������D��   ��EPQQ�$��  �E�� ����E�U���=����}3���G�W��3�����AuB�E���������f�E��E;�})+ȋE��E�t��uG���E��E�t   ��E��m�Iu��E��t���E��3�G��_tj�X  Y�����t�E tj �B  Y���3���^��[��]�U��=|� u%�u�E���T$���\$�$�uj�W  ��$]��$���h��  �u� !   �  �EYY]�U��j �u�u�u�u�u�u�   ��]�U��E3�S3�C�H�EW�  ��H�E�H�M��t�E��  �	X��t�E��  ��H��t�E��  ��H��t�E��  ��H��t�E��  ��H�MV�u�����3A��1A�M����3A��1A�M�����3A��1A�M�����3A��1A��M����3A#�1A�;  ����t�M�I��t�E�H��t�E�H��t�E�H�� t�E	X��   #�t5=   t"=   t;�u)�E��!�M���������M��������E� ���   #�t =   t;�u"�E� ���M�������M�������E�M��3���� 1�E	X �}  t,�E�` �E� �E�X�E	X`�E�]�``�E��XP�:�M�A �����A �E� �E�X�E	X`�M�]�A`�����A`�E��XP�b  �EPjj W�Ȱ�M�At�&��At�&��At�&��At�&��At�&ߋ��������� t/HtHtHu(�   � �%����   ���%����   ��!������� tHtHu!��#�   �	�#�   ��}  ^t�AP���AP�_[]�U��E��t�����w��|��� "   ]���|��� !   ]�U��U�� 3ɋ�9ŀ�t@��|���ń��M��tU�E�E�E�E�E�E��EV�u�E�E h��  �u(�E��E$�u��E��  �E�P�Y������uV�Y���Y�E�^�h��  �u(��  �u�=����E ����]�U���E������W��Dz	��3��   Vf�u�Ʃ�  u|�M�U���� u��tj�ٿ�������Au3�@�3��EuɉM��y���M�O�Et�f�u�U���  f#�f�u��t� �  f�f�u�Ej QQ�$�1   ���#j Q��Q�$�   ���������  ���  ^�E�8_]�U��QQ�M�E�E�����  %�  ���]��f�M��E���]�U��}  ��Eu��u@]Á}  ��u	��ujX]ËM��  f#�f;�uj���  f;�u�E�� u��tj��3�]�jhP������=H�|[�E�@tJ�=�� tA�e� �U�.�E� �8  �t�8  �t3��3�@Ëe�%�� �e��U�E������
�࿉E�U�Ͱ���U��Q�}����E���]�U��Q��}��M�E��#Ef#M�f����E�m�E���]�U��QQ�M��t
�-���]���t����-���]�������t
�-���]����t	�������؛�� t���]����]�U��Q��}��E���]�U��V�u��t�U��t	�M��u��y��j^�0��j����^]�W��+���A��tJu�_��u��ty��j"��3���U��V�u�<��� uV�q   Y��uj褠��Y�4������^]�VW�����S���t�tS�H�S�^���' Y����Ю|�[�> t�~u�6�H�����Ю|�_^�jhp�������=�� u����j�i���h�   ����YY�}3�9���u\j����Y����u�x���    3��Bj
����Y�]�9���uSh�  V�5������4����V��]��Y�E������	   3�@謮���j
�;   Y�VW������~uj �>��h�  �6�ߩ��������Ю|�3�_@^�U��E�4Ű����]����������������SVW�T$�D$�L$URPQQh Td�5    ��3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�-  �   �C��-  �d�    ��_^[ËL$�A   �   t3�D$�H3��4��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�-  3�3�3�3�3���U��SVWj Rh�TQ�T  _^[]�U�l$RQ�t$������]� U����u�M��Si���M��yt~�E�Pj�u��,  ��������   �E�A���}� t�E��`p�����]�U��=�� u�M�P��H��]�j �u����YY]�U����M�SW�u��h���]�   ;�s`�M�yt~�E�PjS�D,  �M������   �X����t�}� ���   �t�E��`p�����   �}� t�M��ap����   �E�xt~-�ÍM����EQ��P�����YY��t�Ej�E��]��E� Y��Uu��3�A� *   �]��E� �E�U�j�pjRQ�M�QW���   �E�P�6(  ��$��u8E��{����E��`p��o�����u�}� �E�t%�M��ap���U��E���Ѐ}� t�M��ap���_[��]�U��=�� u�M�A���w�� ��]�j �u����YY]���WV�t$�L$�|$�����;�v;��h  �%L�s��  ���   ��  ��3Ʃ   u�%����  �%L� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����Z����   u������r*��$�Z��Ǻ   ��r����$�Y�$�Z��$��Y�,YXY|Y#ъ��F�G�F���G������r���$�Z�I #ъ��F���G������r���$�Z�#ъ���������r���$�Z�I �Y�Y�Y�Y�Y�Y�Y�Y�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�Z��Z Z,Z@Z�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$��[�����$�T[�I �Ǻ   ��r��+��$��Z�$��[��Z�Z[�F#шG��������r�����$��[�I �F#шG�F���G������r�����$��[��F#шG�F�G�F���G�������V�������$��[�I X[`[h[p[x[�[�[�[�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��[���[�[�[�[�D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y�����������������U��W�=H���   �}ww�U�����fn��p� ۹   #σ����+�3��of��ft�ft�f��#�uf��#���ǅ�EЃ������Sf��#���3�+�#�I#�[��ǅ�D�_���U��t93���   t�;�Dǅ�t G��   u�fn�f:cG�@�L�B�u�_�ø����#�f��ft �   #Ϻ������f��#�uf��ft@��f����t����뽋}3�������ك��E���8t3�����_��U��UV�uW�z��u� m��j^�0�D^�����   �} v�M� ��~���3�@9Ew	��l��j"���0S�^�Å�~���t��G�j0Z�@I���U�  ��x�?5|�� 0H�89t�� �>1u�B�S�<���@PSV�������3�[_^]�U���,��3ŉE��E�M�SV�uW�u�E�E�E��_���E�3�PWWWWV�E�P�E�P�r.  �؃� �E��t�M��u�E�P��(  YY��u��t��uj���u���tj_�}� t�M܃ap��M���_^3�[�(����]�U���(��3ŉE�SV�u�M�W�u�}�w^���E�3�PSSSSV�E�P�E�P��-  �E�E�WP��"  �ȃ�(�E�u��t��uj�
�u��tj[�}� t�M��ap��M���_^3�[�(����]�U��j �u�u�u������]�U��QQ�ESVW�x�   ��P�ϋ �� �  ������ ���  �}���E���t���  t�� <  �%��  �!��u��u�E!P!f�x�X��<  3����M�����������E�]�s���x&�����ʁ���  ����y�}�}��E�s�f�{_^[��]�U���0��3ŉE��ES�]V�E܍EWP�E�P����YY�E�Pj j���uЋ���f��	4  �u܉C�E��E��C�E�P�uV�0�����$��u�M���_�s3�^[�&����]�3�PPPPP�&[������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��U��M�E������#�V�u�����t$��tj j �=  YY��h��j^�0��Y�����Q�u��t	��<  ����<  YY3�^]�j趏��Y������������U��E3�SVW�H<��A�Y�����t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h��h�d�    P��SVW��1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�jh���#����3����@x��t�e� ���3�@Ëe��E������{V���had� �����U��E���]�U���V�u�M��Y���E�M���E�L0u3�9Ut�E����   �p#E���t3�B�}� ^t�M��ap���]�U��jj �uj ������]�U��} u�u��K��Y]�V�u��u�u�K��Y3��MS�0��uFV�uj �5���԰�؅�u^9��t@V�
���Y��t���v�V�����Y��e���    3�[^]���e������P��e��Y����e������P�e��Y�����U��V�u��tj�3�X��;Es�e���    3��Q�u��uF3Ƀ��wVj�5�����ȅ�u*�=�� tV�\���Y��uЋE��t�봋E��t�    ��^]�U��VW�}��t�M��t�U��u3�f��e��j^�0�FV����_^]Ë�f�> t��Iu��t�+��f��Rf��tIu�3���u�f��d��j"�U��V�u��t�U��t�M��u3�f��d��j^�0��U����^]�W��+��f��If��tJu�3�_��u�f��bd��j"��U��Ef���f��u�+E��H]�U��U�MV��u��u9Mu&3��3��t�E��t��u3�f���u��u3�f��d��j^�0�GU����^]�S��W�����u+��f�3�vf��t%Ou�� +��f��[f��tOtJu��u3�f���_[�{������u�E3�jPf�TA�X�3�f��c��j"�U��E��x!��~��u������������]��Wc���    �T�����]�U���$��3ŉE��ES� �VW�E�3��EV�E��Ӌ��}��
����E�95����   h   Vh�?�а����u&����W�j  VVh�?�а�����S  h�?W�0����?  P��h�?W����0�P��h�?W����0�P��h�?W����0�P�ӣ����th@W�0�P�ӣ���}�� ���t�E��tP�ذ9u�tjX�   9u�t�5����j������;�tO9=��tGP���5���E��ӋM�E��t/��t+�х�t�M�Qj�M�QjP�U��t�E�u�}��    �0���;�t$P�Ӆ�t�Ћ���t���;�tP�Ӆ�tV�Ћ��}�5���Ӆ�tW�u��u�V���3��M�_^3�[�B����]����U�������$�~$�   ��fD$f%�Wf�WfW�f�W��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU@OfV�f($�@@���X��\��Y��Y��Y����X��^�f=�Wf-xW�\�fs�?��fs�?�Y�fp�Df5�W�Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT=pWfs���f%�W���\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<�@O�Y�f(@W�Y��Y��\��X��\��X�f-xW�\��X�f�W�^�f�Wf\�@@���Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5�Wf�f(�Wf(%�WfY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=`Wfp�DfT`W��f%�W���\��Y��X��Y��\����Y��Y��\��\��X��\�f(�Wfp���\��X�fp���X��Y��X�fp���^�f(�Wf(-�Wf(�WfY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(@W�Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$��c��fD$����fD$�D$���f�Wf@WfHW�X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$�������������������U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(Xf(pXf(% Xf(50XfT�fV�fX�f�� %�  f(��Xf(� ]fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(�Xf(�f(�XfY�fY�fX�f(�X�Y�f(-@XfY�f(�PXfT�fX�fX�fY��Y�fX�f(�f�fY˃�f(�f��X��X��X�fD$�D$���fD$f(�X��� f�� �� wH���t^���  wlfD$f(Xf(pXfT�fV���� f�� �� t��Xú�  �OfpX�^�f�X�   �4f�X�Y�������/��������  ���  s:fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$��`���D$���fT$fD$f~�fs� f~с��� ��� t���  릍d$ Q�L$+ȃ����Y�J  Q�L$+ȃ����Y�4  jhИ�H���3��}�j����Y!}�j^�u�;5��}S�������tD�@�tP�j1  Y���tG�}��|)������� P�H�����4��0>��Y����$� F��E������   ���	���Ë}�j����Y�U��V�u��u	V�   Y�/V�,   Y��t�����F @  tV����P�M1  ��YY��3�^]�U��SV�u3ۋF$<uB�F  t9W�>+~��~.W�vV�ś��YP�6�����;�u�F��y����F��N ���_�N�Ãf �^[]�j�   Y�jh������3��}�!}�j�[���Y!}�3��]�u�;5����   �������t]�@�tWPV襚��YY�E�   ������@�t0��uP�����Y���tG�}����u�@tP�����Y���u	E܃e� �   F녋]�}�u����4�V襚��YY��E������   ����t�E��u���Ë]�}�j�����Y�jh������}����������4���3�9^u1j
�a���Y�]�9^uSh�  �FP�~������F�E������*   ���������������P���3�@����Ë}j
�p���Y�U��EVW��x`;��sX���������������Dt=�<�t7�=��u3�+�tHtHuQj��Qj��Qj��ܰ������3����U��� 	   ��U���  ���_^]�U��M���u�U���  ��U��� 	   �B��x&;��s�������������Dt�]��gU���  �U��� 	   ��F�����]�U��M���������������P���]�U���SV�u��t�]��t�> u�E��t3�f�3�^[��]�W�u�M���G���E����    u�M��t�f�3�G�   �E�P�P�e���YY��t@�}��t~';_t|%3�9E��P�u�wtVj	�w�4��}���u;_tr.�~ t(�t�13�9E��3�P�u�E�GWVj	�p�4���u�T������ *   �}� t�M��ap���_�4���U��j �u�u�u�������]�U��Q������u
�..  ������u���  �j �M�Qj�MQP����t�f�E��]����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U��V�u����   �F;�tP�!9��Y�F;�tP�9��Y�F;�tP��8��Y�F;�tP��8��Y�F;��tP��8��Y�F ;��tP��8��Y�F$;��tP�8��Y�F8;�tP�8��Y�F<;�tP�8��Y�F@;�tP�8��Y�FD;�tP�m8��Y�FH; �tP�[8��Y�FL;$�tP�I8��Y^]�U��V�u��tY�;خtP�*8��Y�F;ܮtP�8��Y�F;�tP�8��Y�F0;�tP��7��Y�F4;�tP��7��Y^]�U��V�u���n  �v��7���v�7���v�7���v�7���v�7���v�7���6�7���v �7���v$�7���v(�7���v,�x7���v0�p7���v4�h7���v�`7���v8�X7���v<�P7����@�v@�E7���vD�=7���vH�57���vL�-7���vP�%7���vT�7���vX�7���v\�7���v`�7���vd��6���vh��6���vl��6���vp��6���vt��6���vx��6���v|��6����@���   �6�����   �6�����   �6�����   �6�����   �6�����   �6�����   �}6�����   �r6�����   �g6�����   �\6�����   �Q6�����   �F6�����   �;6�����   �06�����   �%6�����   �6����@���   �6�����   �6�����   ��5�����   ��5�����   ��5�����   ��5�����   ��5�����   �5�����   �5�����   �5�����   �5�����   �5�����   �5�����   �}5����   �r5����  �g5����@��  �Y5����  �N5����  �C5����  �85����  �-5����  �"5����   �5����$  �5����(  �5����,  ��4����0  ��4����4  ��4����8  ��4����<  ��4����@  �4����D  �4����@��H  �4����L  �4����P  �4����T  �4����X  �z4����\  �o4����`  �d4����^]�U��QQ��3ŉE�SV�uW��~!�E��I�8 t@��u������+�H;ƍp|���M$3���u�E� �@�ȉE$3�9E(j j V�u����   PQ�4��ȉM���u3��q  ~Wj�3�X���rKɍA;�v?�E��E   =   w������܅�t���  �P��3����Y��t	���  ���M���M�3ۅ�t�QSV�uj�u$�4�����   �u�j j VS�u�u�S�����������   �E   t,�M ����   ;���   Q�uVS�u�u�������   ��~Oj�3�X����rC�?�A;�v9�}   =   w�������tg���  �P�3����Y��tR���  ���3���tA�E�WVPS�u�u覎������t!3�PP9E uPP��u �uWVP�u$�8���V����YS�ۍ��Y�Ǎe�_^[�M�3���	����]�U����u�M��?���u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap���]�U��Q��3ŉE��MSVW3���u�E� �@�ȉEW3�9E W�u���u��   PQ�4��؅�u3��   ~K�����wC��A;�v9�]   =   w��������t����  �P�1����Y��t����  �������t��PWV�g-����SV�u�uj�u�4���t�uPV�u����V蝌��Y�Ǎe�_^[�M�3������]�U����u�M��u>���u �E��u�u�u�u�uP��������}� t�M��ap���]�U��f�M��  f��f#�f;�u-�EQQ�$����YYHtHtHt3�@]�j�jX]ø   ]��Ɂ� �  f��u�E�� u�} t��Ƀᐍ��   ]��E��������Dz��Ƀ���A@]���Ɂ������   ]�����U��SVWUj j h���u�(  ]_^[��]ËL$�A   �   t2�D$�H�3��k��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    ��3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ�@��SQ�@��L$�K�C�kUQPXY]Y[� ���U����M�S�u�]<���]�C=   w�E苀�   �X�n�ÍM����EQ��P�Ţ��YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�E�PQ�E�P�E�jP�h�������u8E�t�E��`p�3���E�#E�}� t�M��ap�[��]�jh8���~�����95��t*j�Z���Y�e� Vh������YY����E������   ����j����Y�U���D��3ŉE��MSVW�A
3ۋ}��% �  �}��E����  �A���?  �E��A�E�����U��E������u%���9\��u@��|��  3��}𫫫j[�  �\��u��}�UܥH�E�j�]ԥ�H����^#�����Uā�  �yI���A+�3�@�uЋ΃����j^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+ȉ]�3�@���EȋD���M�ȉM�;ȋE؋�j�_r;E�s3�A�MԉD��Jx.��t'�D���ˉ]ԍx;��}؋�r��s3�A�MԉD��JyՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA�X���+\�;�}3��}𫫫������;��  +U܍u�UЍ}��¥��������EċEХ%  �yH���@�EЃ���ǉ]��}Ћ�����j �E�X+�j�E�^�T���ϋ���U�#E؋M����T��C�E�;�|ߋEčU���3�j+Ѓ���E�Y;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��E�3��M�@���D����   �����ЅD���9\��uB;�|��v�}̋�j�Y#������  �yO���G�D��+�3�G��ˉ}���}�;��E�j�_r;E�s3�A�D��Jx(��t!�D���ˍx;��}���r��s3�A�D��Jyۃ���MЋUԋ���!D��B;�}�}��΍<�+�3�����`�A���������E؁�  �yI���A�M܋���j �]��׋]�Y+ˉẺM܋T���ˋ���M�#�U��T���M����E��E�@�E�;�|׋u؍U�����j+�3�Y;�|��D����\����Iy������;T���   �`��}�3�������M�   ��������É�  �yI���A����M�j ��X+��]��׉E؋T������#�U��M����MȉT��C�E�;�|ߋu̍U�����j+�3�Y;�|��D����\����Iy�5h�3�5T�C�   �5h��e�����`�������u�����E؁�  �yI���Aj �]������X+ÉM��׉E܋T���ˋ���U�#ǋM����T��F�E���|ߋ}؍U��uȋ���j+�3�Y;�|��D����\����Iy�}�jX+`��ȋE������%   ��d�u���@u
�E�w���� u�7�M���_^3�[� ����]�U���D��3ŉE��MSVW�A
3ۋ}��% �  �}��E����  �A���?  �E��A�E�����U��E������u%���9\��u@��|��  3��}𫫫j[�  �t��u��}�UܥH�E�j�]ԥ�H����^#�����Uā�  �yI���A+�3�@�uЋ΃����j^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+ȉ]�3�@���EȋD���M�ȉM�;ȋE؋�j�_r;E�s3�A�MԉD��Jx.��t'�D���ˉ]ԍx;��}؋�r��s3�A�MԉD��JyՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA�p���+t�;�}3��}𫫫������;��  +U܍u�UЍ}��¥��������EċEХ%  �yH���@�EЃ���ǉ]��}Ћ�����j �E�X+�j�E�^�T���ϋ���U�#E؋M����T��C�E�;�|ߋEčU���3�j+Ѓ���E�Y;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��E�3��M�@���D����   �����ЅD���9\��uB;�|��v�}̋�j�Y#������  �yO���G�D��+�3�G��ˉ}���}�;��E�j�_r;E�s3�A�D��Jx(��t!�D���ˍx;��}���r��s3�A�D��Jyۃ���MЋUԋ���!D��B;�}�}��΍<�+�3�����x�A���������E؁�  �yI���A�M܋���j �]��׋]�Y+ˉẺM܋T���ˋ���M�#�U��T���M����E��E�@�E�;�|׋u؍U�����j+�3�Y;�|��D����\����Iy������;l���   �x��}�3�������M�   ��������É�  �yI���A����M�j ��X+��]��׉E؋T������#�U��M����MȉT��C�E�;�|ߋu̍U�����j+�3�Y;�|��D����\����Iy�5��3�5l�C�   �5���e�����x�������u�����E؁�  �yI���Aj �]������X+ÉM��׉E܋T���ˋ���U�#ǋM����T��F�E���|ߋ}؍U��uȋ���j+�3�Y;�|��D����\����Iy�}�jX+x��ȋE������%   ��|�u���@u
�E�w���� u�7�M���_^3�[������]�U���   ��3ŉE��E�E��E�E�3�S3�@V�E���É]�W�}��]��]��]��]��]�9E$u�c=���    �.��3��  �U�ʉM��
�� t��	t
��
t��uB��
B�M����{  �$�6��A�<wjXJ�݋E$� ���   � :ujX������+tHHt����  3�@�j� �  X�M��jX�]��3�@�E��A�<v��E$� ���   � :uj묀�+t+��-t&��0t���C�:  ��E~��d���)  j�|���Jj�t����A�<�P����E$� ���   � :�R�����0�c����U���  3�@�E���0|*�E��u���9��s	��0@�G�F�
B��0}�u���E��E$� ���   � :�I�����+�t�����-�k����E���3�@�E��E��E���u��0u�E��
HB��0t��E��E���0|%�u���9��s��0@�GN�
B��0}�u���E���+������-������C~��E�������d�������J�	  3���0@�E���	����j�/����B��E��A�<wj	��������+t"HHt�������j����j���X�M������j����3�@�E���
B��0t���1����   몍A�<v���0�9] t"�B��E�����+t�HH�q����M��jX�z���j
XJ��
�m����H3���@�E����93k�
�u������P  �
B�M���0}���M��Q  ���9�
B��0}�J�E��M���M�����  ��v�E�<|���E��M�OjAX�M���M�����  O8u
HAO8t��M��M�QP�E�P�
  �M�����y��u��E���uu�E���u+u��P  �J  �������/  �����`���  y
���ރ�`9]��  3�f�E���  �ƃ�T���U��u�����  k�� �  ʉM�f9r��}��M��M�����M��y
�U΋�3]�% �  �]ԉE���  #Љ]�#��]܍���  �u�f;��I  f;��@  ���  f;��2  ��?  f;�w�]��7  f��u$F�E�����u�u�}� u�}� u3�f�E��  f��uF�A����u�u	9Yu9t�j�ÍU�_�E��}��}���~X�uč4F�A�E���E��E��M��]�� �ȉM�J�;J�r;M�s3�@��E��J���tf��m���O����M��}��E���@O�E��}�����u��U܁��  �}ԉU�f��~;��x2�E؋�����������U��E�Ҹ��  �}����U��U�f���f��i���  �f��y]�]��������E���E�tC�M؋����M��m�	E��E���������M��U܉E؉}�u�j �ۉU�[tf��3�Gf�f�Eԋ}��f�EԺ �  f;�w���� �� � u@�Eփ��u4�Eډ]փ��u f�E޹��  �]�f;�uf�U�F�f@f�E��@�EڋM��@�E֋M��U���  f;�r3��]�f9E��]���H%   � ���E��:f�E�u�f�EċE؉EƉM�f�u�� 3�f9E���H%   � ���Ẻ]ȉ]ċU��u��������E��MċUƋu����23��ˋË�Ӎ_�#��  �   �j��ˋË����Ë�j�ˋ�[�}�E�f�G
��f��W�w�M�_^3�[������]�T��� �1����.���s�ӐȐ��U���   ��3ŉE��U3�S�]��  V� �  �]�#��E������uA#��E������E����?�U��E�Wf��t�C-��C �}f��u:����   9}��   3��Kf�� �  f;�����$ �C��f�C0 ��  f;���   �E�   �f��M;�u��t�   @uh�i�Gf�}� t=   �u��u0h�i�;�u%��u!h�i�CjP�H���������  �C�h�i�CjP�'���������  �C3��G  �֋�������3ۉ}濈���`f�u��E�   �H�E���  k�Mi�M  �E��?  ������ȋE�E�3�f�E����؉M��E����/  y�ؿ���`�E����  �u��U�u��}���T�}�����  k�� �  ωM�f9r��}čMĉM�����M��y
� �  �E�}����  1E�%�  !u��E�ǉ}�N���E�f;Ƌu��]��]��]�]��}��X  ��  f9M��M��F  f;}��<  f;}�w�]��E  f��u G�E�����}�u��u��u3�f�E��-  f�}� uG�A����}�u	9Yu9t�j�ÍU�^��|����u��u���~r�u��F�q��x����u��u��M��8����B��]��8;ȉM���r;�s3�A��M��B���tf���x����M�������x���N�M�����M��u���|�����@N��|����u����q����}��E����  �u��E�f��~;��x2�E�֋���������E�E���u�����  ��E��E�f���f��q���  �f��ye�]�����3�����E��}�B�}��U�tG�M�����M��m�	E��E���������M��]��E�u�u�j �]����}�[tf��f�f�E��u��f�E� �  f;�w���� �� � u@�E���u4�E��]���u f�E����  �]�f;�uf�M�G�f@f�E��@�E��M��@�E�M���  f;�s f�E�}�f�E��E�E�u��M�U�f�}��!3�f9E���H%   � ���E��Ӊu��U�u��}��E���������M���U�u��E��?  ��f;���  A�]��M��ȋEڋ�3��]��� �  �]�}���  #ǉ]�#ωE������  �}�f;��@  �E�f;E��3  f;}��)  f;}�w�]��2  f��u G�E�����}�u��u��u3�f�E��  f��uG�E�����}�u�}� u�}� t��ӍM�j�U�X����~X�}��E؍<W�E��}����ЋA��]��<;�r;�s3�@��E��y���tf��}��E������}�N�E�����U��E���BH�U��E�����}��u����  f����   �]��]���x,�E�Ӌ���������E�۸��  �]����u�f��Љ]��U�j [f��~[f�M� �  f;�w���� �� � ��   �E�����   �E��]�����   f�E����  �]�f;�u|� �  Gf�E��|�U���  �f��y���������E��}��}��E�tG�]�Ƌ��������������M��]�U�u�j ���u��}�[�M���3�f��@f�f�M��U��<���f@f�E��@�E��u��@�E��  f;�s f�E�}�f�E��E�E�u�U�u�f�}��3�f9E���H%   � ���E����E�M��E��}f�t6���}���/3�f�� �  f9E�����$ �A3�@�A�A0�Y�  �}�jX;�~�E��}������?  3�j�}�f�E�]�_�ʋ���������Љu��]�Ou�}��]��U�u�j [��y7�߁��   ~-�]����������������O�]�u����]�3ۉU�u��u��E�@�E��~�}��ωM�����   �u��ʍ}����ҥ��}������ЋE��4 ��������������E��8�M�;�r;�s�B��;�r��s3�A�ɋЋM�tF�Eȍ<;�r;�sFű��U�������U��U��?����6�U���M��E���0�]�A�E�H�M��E���~�E�E��>����u��}��A���<5|E�	�99u�0I;�s�;�sAf���E�*Ȁ��H�Ɉ\3�@�M�_^3�[�[�����]À90uI;�s�;�s̋M�3�f�� �  f9E�����$ �A3�@�A�0����3�SSSSS����U��M3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tƋѻ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t;�u �  ]Ã�@]�@�  ]�U�����}�f�E�3ɨtjY�t���t���t��� t���t��   SV��   ��W�   #�t&��   t��   t;�u��   �
����   ��   t;�u��   ���   ���   ��t��   �}���E��#�#��;���   V�?  ��Y�E��m���}��E�3��tj^�t���t���t��� t���t��   �Ћ�#�t*��   t��   t;�u��   ���   ���   ��   t��   u��   ���   �   ��t��   �=H���  ���]�E�3Ʉ�yjY�   t���   t���   t����t���   t��   �л `  #�t*��    t�� @  t;�u��   ���   ���   j@%@�  [+�t-�  t+�u��   ���   ���   ��#}��#��;���   P�$���P�E�t���YY�]�E3Ʉ�yjY�   t���   t���   t���   t���   t��   �п `  #�t*��    t�� @  t;�u��   ���   ���   %@�  +�t-�  t+�u��   ���   ���   ���3Ʃ t��   ������_^[��]�U��M3���t@��t����t����t����t�� ��   t��V�Ѿ   W�   #�t#��   t;�t;�u   �   �   �с�   t��   u���_^��   t   ]�U��V�uW�����u��'���    �!����E�F�t9V�t���V���   V�[k��P�  ����y�����~ t�v����f Y�f ��_^]�jhX��]������}�3��u������u�a'���    ������]����F@t�f ��V�j��Y�e� V�?���Y���}��E������   �ǋu�}�V�Pj��Y�jhx��%]��3��u�}���u��&��� 	   �   ����   ;=����   �����E��߃��������D��trW����Y�u��E������Dt(W����YP����u�����u��t�<&���0�i&��� 	   ����u��E������
   ���!�}�u�W����Y��:&��� 	   �}������\��á�����t���tP���3�PPjPjh   @h�i������U���S�]3ҸN@  VW�E���S�S9U�<  �ʉU�M�U��U�}�����ҥ���u�΋}��������������������E����s{3ɉE;�r;E�s3�A���t��3ɍp;�r��s3�A�s��tG�{�U�3���M�;�r;�s3�@�K��tG�{�U�u��}���e� �������E���s�{� �u�}��E��M�;�r;�s3�@��E����t$��3ҍp�u;�r��s3�B�s��tG�}��{�EH�s�E�{�E��������N@  3�9Su.�S������������E�����  ��E���tۉS�s�S�� �  u4�;�s�ǋ��������E�����  ��E��� �  tى;�s�S_^f�C
[��]�jh���&Z��3ۉ]�u���u�#�����#��� 	   �   ����   ;5��s{���������������D8��u
�y#���  �ZV����Y�e� �����D8tV�T   Y����#��� 	   ����}��E������
   ���(�u�}�V�����Y��#����I#��� 	   �������Y���U��VW�}W�=���Y���tP�����u	���   u��u�@Dtj����j���	���YY;�tW�����YP����u
�����3�W�Y���Y�σ����������D9 ��tV�"��Y����3�_^]�U��V�u�F�t �Ft�v�����f����3�Y��F�F^]�������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �������������%��%̰���̃=�� uK�x���t���Q�@<�@�Ѓ��x�    V�5����t������V���������    ^�                                                                           ,� <� L� ^� t� �� �� �� �� ̛ ܛ �  � � (� >� P� `� n� �� �� �� Ȝ ޜ �� � ,� H� f� �� �� �� �� ʝ ؝ � � � � &� 2� B� Z� r� �� �� �� �� Ğ О ܞ � �� � � 0� @� P� b� v� ��                   ��J�Z���        ��H�                    ߃DT       O   j X     ߃DT          hj hX                      ������������       ����       ����       ����                     ������������       ����       ����       ����         ����    ����������������   ��������       ����   �������� k��  �0�@�P�`�p�����    0   .   -   ||----------------------------------------  ||  (c) 2012-2014 - Christopher Montesano   ||  http://www.cmstuff.com   v  ||      ||    build date:   �l�� ����d ����������� ���`N��gui_icons.tif   gui res mp� �� p�@p� `p`@��?�?`�?�?�?0�@b��p@�@�@ �   %  `m��  dp� P`���@�e:\repos\cmnodes\src\source\customgui\cmcustomguireal.h CM_REAL_GUI cmRealGUI   �m�� ���������������� �� �0�@�P�`�p� ���e:\repos\cmnodes\src\source\prefsdialog\cm_prefs.h  Prefs_cm    cmStuff @n�� ���������������� ��0��@���`�p�`���e:\repos\cmnodes\src\source\prefsdialog\cmnodes_prefs.h �n� Є�������������� �� �0�@�P�`�p�e:\repos\cmnodes\src\source\nodes\cmnodetree.h  �nЧ `� P��`�p� � �����P� �0�@�P�`�p��������  0cmNodeTreeRoot  cmNodeBaseRoot  0123456789  StartUndo 11    AddUndo 13  EndUndo 11  AddUndo 14  AddUndo 15  AddUndo 16  AddUndo 17  AddUndo 18  AddUndo 19  e:\repos\cmnodes\src\source\scenehook\cmnodeforest.h    8o� �a@c�����c�e���� �� �0�`cPc`�p�@� 4`� h����0n�ip�Pme:\repos\cmnodes\src\source\nodes\node_types\cmnodeoutput.h input   �o � ��@c�������e���� �� �0�`cPc`�p�@� N`� h����l�i i�~�d�AAddUndo 20  AddUndo 21  StartUndo 14    EndUndo 14  color   diffusion   luminance   transparency    reflection  environment bump    normal  alpha   specular    displacement    p`�  �@c�����c�e���� �� �0�`cPc`�p��Ip��ep���@n�i��Pme:\repos\cmnodes\src\source\nodes\node_types\cmnodeinput.h  pp��  �@c�����c�e���� �� �0�`cPc`�p���`��ep���@n�i��Pm�pЪ 0�@c�����c�e���� �� �0�`cPc`�p����A`� ep�0�pl�ip�Pme:\repos\cmnodes\src\source\nodes\node_types\cmnodechannels.h   q�� ��@c�����c�e���� �� �0��]Pc`�p�p��`� ep��}k�i�hPminputA  inputB  lq � ��@c�����c�e���� �� �0�`c0�`�p�0� �`� ep���@k�iiPmNormal  Darken  Multiply    Color Burn  Linear Burn Darker Color    Lighten Screen  Color Dodge Linear Dodge    Lighter Color   Overlay Soft Light  Hard Light  Vivid Light Linear Light    Pin Light   Hard Mix    Difference  Exclusion   Subtract    Divide  Hue Saturation  Color   Luminosity  Levr    Grain Extract   Grain Merge mask    �qP� ��@c�����c�e���� �� �0�`c��`�p�P�&`�@fp���@k�iiPme:\repos\cmnodes\src\source\nodes\node_types\cmnodeadjust.h Add Minimum Maximum r`� @�@c�����c�e���� �� �0�]Pc`�p��p�`�@fp��}l�i�hPmhr�� @�@c�����c�e���� �� �0�`cPc`�p�P���`�@fp��}l�i�hPm�r`�  �@c�����c�e���� �� �0�`cPc`�p����`�@fp��}l�i�hPms0� ��@c�����c�e���� �� �0�`c`�`�p�0�0�`�@fp�0�pl�ip�PmLinear -> Linear    Linear  HSV HSL sRGB     ->     ds��  �@c�����c�e���� �� �0��^Pc`�p�p�`�@fp��}l�i�hPm�s� `�@c�����c�e���� �� �0�`cPc`�p���P�0�@fp���pl�ip�Pmt� p�@c�����c�e���� �� �0�`cPc`�p�@�0$`�@fp��}l�i�hPm`t�  �@c�����c�e���� �� �0�`cPc`�p���PL`��gp�0�pl�ip�Pme:\repos\cmnodes\src\source\nodes\node_types\cmnodeeffects.h    �t�� �@c�����c�e���� �� �0�`cPc`�p� �`��gp� @k�iiPmsource  displace    up� P�@c�����c�e���� �� �0�`cPc`�p����`��gp��}l�i�hPm\u�� ��@c�����c�e���� �� �0�`cPc`�p����*`��gp��}l�i�hPm�u0� `�@c�����c�e���� �� �0�\Pc`�p�����`��gp��}l�i�hPmv�� �@c�����c�e���� �� �0�`cPc`�p� ��`��gp���pl�ip�PmXv � У@c�����c�e���� �� �0� ^Pc`�p� ��`��gp��}l�i�hPm�v�� Ъ@c�����c�e���� �� �0� _Pc`�p��� `��gp���pl�ip�Pm w�� P�@c�������e���� �� �0��_P�`�p�`�P`��fp���@n�i��PmFacing Ratio    UV Coordinates  Camera Distance Normals (Object)    Normals (World) Normals (Camera)    Object Color    Normal Direction    e:\repos\cmnodes\src\source\nodes\node_types\cmnodeutility.h    Tw � ��@c�����c�e���� �� �0�`cPc`�p�@� C`��fp��~pl�ip�Pm�wP� ��@c�����c�e���� �� �0�`cPc`�p� �@ `��fp��~@n�i��Pm�w0� p�@c�����c�e���� �� �0�`c��`�p����H`��fp�ЁPn@j iPminput 0 input   Pxp� p�@c�������e���� �� �0��aPc`�p����9`��fp���@n�i��Pm�x�� �a@c�����c�e���� �� �0�`cPc`�p�@�/`��fp�0�pljp�Pm�x�  �@c�����c�e���� �� �0�`cPc`�p����`��fp�`~pl�ip�PmLy0� ��@c�����c�e���� �� �0�`cPc`�p�� `��fp���@n�i��Pm�y�� �a@c�����c�e���� �� �0�`cPc`�p�@��I`��fp���n�j0iPmtile    �y�� ��@c�����c�e���� �� �0�`cPc`�p�p�P?`��fp���@n�i��PmHz� P�@c�����c�e���� �� �0�`cPc`�p����/`��fp���pl�ip�Pm�z`� ��@c�����c�e���� �� �0�`cPc`�p�����`��fp��|�jPi iPmcontrol �z@� �@c�����c�e���� �� �0� aPc`�p�`��4`��fp���pl�ip�PmD{@� p�@c�������e���� ��pT0�`cPc`�p�@� N`��h�����n�i@i�~�d�BAddUndo 22  AddUndo 23  StartUndo 15    EndUndo 15  e:\repos\cmnodes\src\source\nodes\node_types\cmnodevray.h   matte opacity   matte alpha material weight luminosity color    luminosity dirt luminosity occulded luminosity unocculded   luminosity transparency flakes color    flakes glossiness   flakes orientation  reflection color    reflection transparency specular1 color specular1 transparency  specular1 hilight glossiness    specular1 reflection glossiness specular1 anisotropy    specular1 anisotropy rotation   specular1 reflectance 90 degree specular1 reflectance 0 degree  specular2 color specular2 transparency  specular2 hilight glossiness    specular2 reflection glossiness specular2 anisotropy    specular2 anisotropy rotation   specular2 reflectance 90 degree specular2 reflectance 0 degree  specular3 color specular3 transparency  specular3 hilight glossiness    specular3 reflection glossiness specular3 anisotropy    specular3 anisotropy rotation   specular3 reflectance 90 degree specular3 reflectance 0 degree  specular4 color specular4 transparency  specular4 hilight glossiness    specular4 reflection glossiness specular4 anisotropy    specular4 anisotropy rotation   specular4 reflectance 90 degree specular4 reflectance 0 degree  specular5 color specular5 transparency  specular5 hilight glossiness    specular5 reflection glossiness specular5 anisotropy    specular5 anisotropy rotation   specular5 reflectance 90 degree specular5 reflectance 0 degree  diffuse1 color  diffuse1 dirt   diffuse1 occulded   diffuse1 unocculded diffuse1 transparency   diffuse1 roughness  diffuse2 color  diffuse2 dirt   diffuse2 occulded   diffuse2 unocculded diffuse2 transparency   diffuse2 roughness  refraction color    refraction glossiness   refraction translucency sss overall color   sss color   sss scatter color   sss scatter radius  AddUndo 2   �{��  D0�@�p�`�p�����e:\repos\cmnodes\src\source\command\cmnode_commands.h   cut.tif #$  �{�� �C0�@�p�`�p�����copy.tif    8|�� �D0�@�p�`�p�����paste.tif   �|��  D0�@�p�`�p�����delete.tif  �|��  E0�@�p�`�p�����select_all.tif  (}�� @D0�@�p�`�p�����deselect_all.tif    x}�� `D0�@�p�`�p�����disconnect.tif  �}�� �D0�@�p�`�p�����frame_selected.tif  ~�� �D0�@�p�`�p�����preferences.tif h~�� �C0�@�p�`�p�����add_tree.tif    �~�� @E0�@�p�`�p�����tree_menu.tif   �� �D0�@�p�`�p�����node_menu.tif   X�� �E0�@�p�`�p�����zoom_in.tif ��� �E0�@�p�`�p�����zoom_out.tif    ��� `E0�@�p�`�p�����zoom_100.tif    H���  E0�@�p�`�p�����reset_view.tif  ���� �C0�@�p�`�p�����calc_preview.tif    03  04  05  06  #$07--  08  09  10  11  #$12--  13  #$14--  15  16  17  #$18--  19  20  21  22  23  ��� �I0�@�p�`�p����� node   Create  node_solid_color.tif    8���  J0�@�p�`�p�����node_texture.tif    ����  F0�@�p�`�p�����node_clamp.tif  ؁�� @F0�@�p�`�p�����node_colorspace.tif (��� �F0�@�p�`�p�����node_curves.tif x��� �G0�@�p�`�p�����node_filter.tif Ȃ�� �G0�@�p�`�p�����node_grade.tif  ��� �H0�@�p�`�p�����node_math.tif   h��� �E0�@�p�`�p�����node_blend.tif  ���� �F0�@�p�`�p�����node_copy.tif   ��� �I0�@�p�`�p�����node_shuffle.tif    X��� �E0�@�p�`�p�����node_blur.tif   ���� �F0�@�p�`�p�����node_dirblur.tif    ����  G0�@�p�`�p�����node_distort.tif    H��� @G0�@�p�`�p�����node_edge_detect.tif    ���� `G0�@�p�`�p�����node_emboss.tif ��� �H0�@�p�`�p�����node_matrix.tif 8��� �H0�@�p�`�p�����node_normal_map.tif ���� @J0�@�p�`�p�����node_transform.tif  ؆��  I0�@�p�`�p�����node_output.tif (��� `H0�@�p�`�p�����node_material.tif   x���  F0�@�p�`�p�����node_colorize.tif   ȇ��  H0�@�p�`�p�����node_info.tif   ��� �G0�@�p�`�p�����node_highpass.tif   h��� �I0�@�p�`�p�����node_switch.tif ���� @H0�@�p�`�p�����node_invert.tif ��� �I0�@�p�`�p�����node_specular.tif   X��� `J0�@�p�`�p�����node_vrayadvanced.tif   ����  G0�@�p�`�p�����node_distance.tif   ���� @I0�@�p�`�p�����node_reflection.tif H��� �H0�@�p�`�p�����node_noop.tif   ���� �F0�@�p�`�p�����node_diffuse.tif    ��� �G0�@�p�`�p�����node_fresnel.tif    8���  J0�@�p�`�p�����node_tiler.tif  ���� `I0�@�p�`�p�����node_shadow.tif ؋�� `F0�@�p�`�p�����node_condition.tif  (���  I0�@�p�`�p�����node_projector.tif  x���  H0�@�p�`�p�����node_input.tif  ?   Are you sure you want to delete bookmark     has been saved.    Bookmark    ��� �J0�@���`�p�����Tree Bookmark 01    e:\repos\cmnodes\src\source\command\cmtree_bookmark_commands.h  tree_bookmark.tif   X��� �J0�@���`�p�����Tree Bookmark 02    ���� �J0�@���`�p�����Tree Bookmark 03     ��� �J0�@���`�p�����Tree Bookmark 04    T��� �J0�@���`�p�����Tree Bookmark 05    ���� �J0�@���`�p�����Tree Bookmark 06    ���� �J0�@���`�p�����Tree Bookmark 07    P��� �J0�@���`�p�����Tree Bookmark 08    ���� �J0�@���`�p�����Tree Bookmark 09    ���� �J0�@���`�p�����Tree Bookmark 10    0,0 %.0f,%.0f   %.2f    L�@� ��0���`���@� �����Cut Copy    Paste   Delete  Disconnect  Calculate Previews  StartUndo 10    AddUndo 3   AddUndo 4   EndUndo 10  New Tree    StartUndo 2 AddUndo 5   AddUndo 6   EndUndo 2   Error: Could not initialize copy operation  AddUndo 7   cmNodeMat   cmNodeVrayAdv   StartUndo 3 AddUndo 8   EndUndo 3   Error: Could not initialize paste operation StartUndo 4 AddUndo 10  AddUndo 11  AddUndo 12  AddUndo 28  EndUndo 4   unknown StartUndo 5 EndUndo 5   StartUndo 6 EndUndo 6   StartUndo 7 EndUndo 7   StartUndo 8 EndUndo 8   No tree selected    StartUndo 9 EndUndo 9   Add Tree... &c& ���  � p��� P`p�� � Edit    View    Nodes   Bookmark    cmNodeEditor    �� �J0�@�p�`������4�� �� �� � P� `���@�File    New...  Load... Save... Save All... Copy All    Delete...   Rename...   load    selection   StartUndo 13    AddUndo 25  AddUndo 26  AddUndo 27  EndUndo 13  Are you sure you want to delete     cmtree  Load    Save    cmTreeManager   ���� �M0�@�p�`������Б � ����0�cmUpdateNodeThread  e:\repos\cmnodes\src\source\utility\cmbghandler.h   P��� `| �������| � ���� �� �0� P�`�p�`p } �~ �~ ����e:\repos\cmnodes\src\source\shader\cmnodeshader.h   Could not find string resource for node     Could not find string resource for category      description    Failed to register  nbase.tif   Node limit exceeded Scmnodeforest   Failed to register cmNodeForest description cmNodes Failed to register cmNodeForest cmNodeTree  Failed to register cmNodeTree   Nbase   Ncolor  Ntexture    Nclamp  Ncolorize   Ncolorspace Ncurves Nfilter Ngrade  Ninvert Nmath   Nblend  Ncopy   Nshuffle    Nblur   Ndirblur    Ndistort    Nedgedetect Nemboss Nhighpass   Nmatrix Ntransform  Noutput Nmaterial   Nvrayadvanced   Ncondition  Ndiffuse    Ndistance   Nfresnel    Ninfo   Nnoop   Nnormalmap  Nprojector  Nreflection Nshadow Nspecular   Nswitch Ntiler  e:\repos\cmnodes\src\source\utility\cmnoderegister.h    #$00cmNodeEditor    Failed to register cmNodeEditor #$01cmTreeManager   Failed to register cmTreeManager    #$02--  cmNode  Failed to register AM Hook  xcmnodeshader   cmNodeShader    prefs_cmnodes   e:\repos\cmnodes\src\source\main.cpp     R13    1001;   1002;   1003;   1004;   1005;   1006;   1007;   Component Failure:  Shaders Cinema4D                ���ư>-C��6?{�G�zt?#���?�������?)\���(�?]m���{�?�������?�v��/�?333333�?
ףp=
�?�������?���z6�?      �?�Q����?���(\��?�A`��"�?333333�?UUUUUU�?�������?]t�E�?      �?�p=
ף�?�(\����?bX9���?333333�?UUUUUU�?�,C���?      �?�������?ffffff�?      �?�z�G��?�������?       @333333@      @      @-DT�!	@      @      @      @-DT�!@       @      "@ףp=
�)@      4@      >@      Y@     �b@     �f@     �o@     @@     @�@������      �      �333333�              �?              �?{�G�zt?�������?�������?�������?�������?333333�?333333�?�(\����?��(\���?�������?�������?      �?      �?��Q���?      �?333333�?333333�?      �?      �?333333�?333333�?���Q��?)\���(�?
ףp=
�?�������?)\���(�?���Q��?      �?      �?�������?�������?ףp=
��?333333�?�G�z��?)\���(�?              �?{�G�zt?      �?�������?      �?      �?      �?      Y@      Y@��������������������������       �       ����������������� }�a@c�����c�e���� �� �0�`cPc`�p�`h j�jk�k�kl l@mPmoutput  CopyTo - Update StartUndo 1 AddUndo 1   EndUndo 1   TRUE    FALSE   SetNodeDirty:            �V@              �?�������?�������?      �?      �?�������?�������?      �?����c:\program files\maxon\cinema 4d r13\resource\_api\c4d_file.cpp c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basebitmap.cpp   ̒0��������W������ ��`������������V 0@P`p����V 0@P`p� 9���V 0@P`p��=h��V 0@P`p� ?�?�?�?�?�?�?�?�?`@p@�@�@c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gui.cpp  ~   Progress Thread 0%  %   ��������h㈵��>����MbP?
ףp=
�?-DT�!�?      �A-DT�!��       �        -DT�!�?              �A        -DT�!��c:\program files\maxon\cinema 4d r13\resource\_api\c4d_general.h       %s  |�0�p���p�c:\program files\maxon\cinema 4d r13\resource\_api\c4d_baseobject.cpp   D���������p�c:\program files\maxon\cinema 4d r13\resource\_api\c4d_resource.cpp #   M_EDITOR    ؔ�� ���������������� �� �0�@�P�`�p� ���    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp    ��S4��S|�pS    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gv\ge_mtools.cpp ĕ@Tc:\program files\maxon\cinema 4d r13\resource\_api\c4d_basetime.cpp        ����A  4&�kC �Ngm��C  4&�k�c:\program files\maxon\cinema 4d r13\resource\_api\c4d_libs\lib_ngon.cpp        fmod         t�&���&���&���&���������&�&���&�      8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7      �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC                                            �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               �       �      ��      ������    ����    ��      ��            8C      8C      0<      0<��+eGW@��+eGW@  ��B.�?  ��B.�?:;����=:;����=�ѱt�?Z�fUUU�?���&WU�?{������?                Mu�{�<`�w>�,  �g5RҌ<t�ӰY  a��aN�`<țuE�  l{�]���<��lX�  ќ/p=�><���2��  ؼcnQ�<P[� {8�&TŤ<�-���B �?RbSQ�<zQ}<�r �S?���<u�o�[� _/:>��<��h1�� �æDAo�<֌b�; �������<8bunz8 ���+G�<�|�eEk 1�	m���<����� �
r�7�<䦅� ���MuM�<�1
� J��]9ݏ<�d�< )}̌/�<ʩ:7�q �^�s)ҧ<���4ۧ mL*�H��<"4L�� ��%F��<).�!
 ��`�cC<-�a`N y����n<�<���� ��z�ΐv<'*6�ڿ 	*(�̃�<�,�v�� ���	�<�O�V+4 ���5�<�'�6Go 	T��c�<)TH�� 5�d+�2�<H!�o� 
���<�U:�~$ �s ��<$"U�8b qU�M��<�;f�� �GΆ�+�<.e<�� �o � �<s_��u ���"a�<�gBV�_ ��F�D�<��s� Ul֫��e<bN�6�� �g�����<�L��% ���<�D��h ����/��<۠*B� D_�Y��{<6w��� <(��`�<��Ͱ77	 �b� ��<ONޟ�}	 'Α+��q<�𣂑�	 �.�X4m�<d�]{f
 ����|'�<\%>�U
 �Zsn�i�<��yUk�
 �3˒w�<��Z���
 �-�f$�<�O��3 ���.�<F^��v ��_
��t<��K�� ��0�ns<�R�ݛ �Y	я��<K�W.�g h�l,kg<i��� � ���6	p�<{�J- �=���t<����X ����PZ�<�2�� ��Js��<^�{3�� ӈ:`�t<�?��.P &I	�'o�<ِ����  �A�Î<'Za�� ��1�d�<@En[vP �͑M;�w<ؐ����       �?       �9��B.�@  ׽2b      �        �������         0<  0<�dW�dW      �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �      �?      �?3      3                      �                     �              �?      �?3      3            �      0C       �       ��              �~���          8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �        ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=(null)  ( n u l l )            EEE50 P    ( 8PX 700WP        `h````  xpxxxx          (�x�    �������             ��      �@      �               ���5�h!����?      �?            �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��log log10   exp pow asin    acos    exp10   atan    ceil    floor   modf    sin cos tan sqrt       �U��?�wB%�K�=      �?   �[��?(�6N�g�=      �?   $�?V�`t� >      �?   ��տ?��2n{a>      �?   ����?��M��=      �?   H{��?{4�r>      �?   Pא�?"�"�>      �?   �u[�?��*��>      �?   ����?G�0��_(>      �?   4wb�?��i^^?(>      �?   ��0�?p3���>      �?   @��?F��M>      �?   8M��?�B�V��>      �?   ��d�?}B��a.>      �?   ȴ�?d�����>      �?   g��?�ߊ��>      �?   �@�?�f\���*>      �?   �~e�?�-��f>      �?   �]%�?D	�G��?>      �?   ���?�\����>>      �?   X���?�1��#>      �?   �E�?��h��>      �?   �?��?�ⳇ��>      �?   ����?�$	�49>      �?   x�8�?k���0H<>      �?   ����?r��ش8>      �?   8fm�?�"m>">      �?   ħ �?[��<c�'>      �?   �k��?"���%>      �?   ���?݉@fR�8>      �?   ����?��T���:>      �?   T�!�?3&�F>      �?   � ��?<����[#>     ��?   �%�?�Y:/(A6>      �?   ����?��N��2>     ��?   8O�?�r�!'	>      �?   ��r�?���8{K>     ��?   �p��?9��l�9$>      �?   �
G�?�aj	�i9>     ��?   T|��?'\�|#<>      �?   $��?�}�dj�#>     ��?   �Wn�?׈MVx:>      �?   ,���?1�8o,>     ��?   D�$�?	c�/�
>      �?   @ |�?��x7|�1>     ��?   |���?��9>      �?   p #�?�IA��u=>     ��?   �s�?�x ٴ4>      �?   p���?edf�&�.>     ��?   ,�?��f���A>      �?   h�*�?v����2>     ��?   $gN�?RE\��K>      �?   �q�?'^��IE>     ��?   DΒ�?��&a��H>      �?   L���?�&KrQF>     ��?   ,���?�#/�'�>      �?   إ��?]X�c�?>     ��?    ��?�Ԯ}�>      �?   �e.�?�IdW�A>     ��?   �K�?���ΐ?>      �?   Xg�?��4*�A>     ��?   _��?�[�ǆJ>      �?   ���?1���0H>     ��?   ���?�hc#�]G>       @   ,*��?�Q�x
�F>     @ @   p���?ek�R�.N>     � @   �� �?�Ӿ�n@>     � @   �b�?�����O>      @   $Q/�?CJ���O>     @@   ��E�?������G>     �@   �[�?�3E�{A>     �@   T�p�?�SfI�S:>      @   X΅�?B6)�1�<>     @@   �3��?>ځ���7>     �@   $��?s(��N>     �@   @���?V�
6�f=>      @   (���?��{��>     @@   (W��?��-�Jg >     �@   ����?��"a�PK>     �@   xm�?,S��ڤ6>      @   ���?�6��hb">     @@    �-�?�k,�<>     �@   X�>�?�0����=>     �@   �O�?�׀IX�H>      @   �-_�?���
@>     @@   ��n�?���2E>     �@   �P~�?�=�ő�8>     �@   lj��?�[j&,>      @   L7��?��x��82>     @@   ����?c�#V�B>     �@   0��?7ڨ.�Y>     �@   P���?�[�p&>      @   ؔ��?h4�M��A>     @@   � ��?E�p�l E>     �@   �+��?�o�$�E>     �@   h��?\���*�K>      @   ���?-�?��B>     @@   P8�?�(l�|�@>     �@   �p!�?u���@�J>     �@   @p-�?�V��1>      	@   �89�?����5>     @	@   <�D�?��ƀ�7>     �	@   h)P�?R`D�OG>     �	@   �T[�?9%� ��K>      
@   �Mf�?��/�<>     @
@   �q�?�Ò��?>     �
@   �{�?4��2G<>     �
@   L��?Â���|/>      @   �Y��?���s�
@>     @@   �k��?��Ò�a@>     �@   XS��?x(3��u8>     �@   ���?v�O,ib>      @   ȥ��?�&L͒C>     @@   ���?��}��L>     �@   �X��?Lo����>     �@   �x��?-�Ϡ�9>      @   �s��?6FID?9>     @@   8J��?����gsL>     �@   d���?��y>     �@   ���?>�&�09C>      @   ����?
��<�A>     @@   (J�?I�V	C>     �@   `w�?��^@�N>     �@   ���?�#��%�@>      @   �s�? �M�K>     @@    D'�?ή�Q��->     �@   ��.�?9!���G>     �@   ��6�?.����1>      @   >�?.1�NcB>      @   �cE�?�sǔ�1>     @@   L�L�?�n�HN>     `@   H�S�?�W��$>     �@   8�Z�?
Ȃ�q�;>     �@   ��a�?N�/�[7>     �@   (�h�?�=�mC>     �@   0oo�?�H75M>      @   Hv�?P��.�#>      @   �|�?�G���7>     @@   �*��?�#4��2I>     `@   ����?o���oJ>     �@   ����?���-��#>     �@   ���?�h��%F>     �@   @��?R�x^D>     �@   PP��?�� s�@>      @   4L��?P�_!
�#>      @   4��?��:#�G>     @@   L��?qg�:&J>     `@   Hɹ�?5L$.��4>     �@   \w��?!�1�C>     �@   ���?���[<>     �@   D���?��<���=     �@   ���?��
~���=      @   �y��?������B>      @   ����?�~.���4>     @@   h��?��u�|�8>     `@   �E��?A8yL;>     �@   �h��?��41��C>     �@   �{��?-���+oF>     �@   $��?x���O>     �@   s��?�՝m�T2>      @   �W��?����=>      @   �-�?î�\�=>     @@   ��?���\=�=     `@   ��?j\&">     �@   �X�?��1�D>>     �@   ���?�#O#`�I>     �@   ��?�}���0>     �@   ��?���F\IE>      @   t{#�?��ׯ,B>      @   0�'�?�E� ]�$>     @@   ,>,�?��ކ?5>     `@   ��0�?��iIqE>     �@   ��4�?�ha�;>     �@   �9�?��A���D>     �@   �.=�?̤KF�w�=     �@   DMA�?�����=      @   `E�?ap�I0�H>      @   �gI�?��:���->     @@   �cM�?��%Q>     `@   @UQ�?Ly5ښoE>     �@   �;U�?v�g�0�/>     �@   �Y�?jv�U�G>     �@   �\�?�����yK>     �@   ,�`�?A%My��>      @   md�?���H>      @    h�?�p���M>     @@   0�k�?k��}<>     `@   �ho�?����f7O>     �@   ��r�?���}�O>     �@    �v�?+��i�I>     �@   @z�?�b�B'=>>     �@   `�}�?Z����M>      @   ����?1�����M>      @   �a��?R�~���=     @@   t���?QNT	��B>     `@   x��?�W3c�L>     �@   g��?�+(����=     �@   D���?q���J�K>     �@   L��?� ;,*>     �@   8!��?������D>      @   ,O��?� ����E>      @   Du��?��in]D>     @@   ����?%����3F>     `@   P���?^��F"VM>     �@   ����?�}�30}->     �@   @���?�~F	y�;>     �@   ����?l	R(>     �@   躰�?��\�7`>      @    ���?�dg���;>      @   ���?�;Sv�@E>     @@   <|��?�����M>     `@   �Y��?|}�;�2>     �@   ,0��?�<v��G>     �@   $ ��?̯�/p�">     �@   ����?���\(0>     �@   |���?[s$���F>      @   I��?�d�ӔV>      @   T���?���0)LK>     @@   h���?�)�5G�5>     `@   XY��?�|��zJ>     �@   @���?W�޾�L?>     �@   0���?����6:>     �@   <3��?��Q���B>     �@   x���?7o��/�M>      @   �Q��?�Kc�Z�0>      @   ����?�z-�A5>     @@   Z��?"B�DcI>     `@   ����?��`I�.>     �@    L��?L�d�%>     �@   ���?"�l"w �=     �@   �(��?�?��!>     �@   ���?��j^�J>      @   8���? ϞH��0>      @   LL��?���%�C>     @@   T���?��J�+N>     `@   d���?;l�>�0>     �@   �B��?�^{v�@>     �@   Ȋ��?�@Y˕B>     �@   @� �?T�l���0>     �@   ��?w4n4>      @    G�?�oN�=�;>      @   h|�?�L�{�/>     @@   <�	�?B�nu5>     `@   ���?���`�,+>     �@   d�?����5>     �@   �$�?l��  >     �@   �C�?~+^��M>     �@   �^�?�PK�QD >      @   ,u�?^{�#tF>      @   |��?�^4K�� >     @@   ���?��4�O
>>     `@   ���?XEړ� J>     �@   ���?(�gԹ�,>     �@   �� �?43-spF>     �@   ��"�?P`E5�+*>     �@   ��$�?=�QQ�D>       @-DT�!�?\3&��<e+000     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          �      	   m s c o r e e . d l l   CorExitProcess  k e r n e l 3 2 . d l l     FlsAlloc    FlsFree FlsGetValue FlsSetValue InitializeCriticalSectionEx CreateEventExW  CreateSemaphoreExW  SetThreadStackGuarantee CreateThreadpoolTimer   SetThreadpoolTimer  WaitForThreadpoolTimerCallbacks CloseThreadpoolTimer    CreateThreadpoolWait    SetThreadpoolWait   CloseThreadpoolWait FlushProcessWriteBuffers    FreeLibraryWhenCallbackReturns  GetCurrentProcessorNumber   GetLogicalProcessorInformation  CreateSymbolicLinkW SetDefaultDllDirectories    EnumSystemLocalesEx CompareStringEx GetDateFormatEx GetLocaleInfoEx GetTimeFormatEx GetUserDefaultLocaleName    IsValidLocaleName   LCMapStringEx   GetCurrentPackageId GetTickCount64  GetFileInformationByHandleExW   SetFileInformationByHandleW    П   0�	   ��
   �   (�   ��   �   (�   ��   �   @�   ��    �   l�   ��    x�!   �"   Чx   8�y   X�z   t��   ���   ��R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
         R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
         R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 4  
 -   i n c o n s i s t e n t   o n e x i t   b e g i n - e n d   v a r i a b l e s  
     D O M A I N   e r r o r  
     S I N G   e r r o r  
     T L O S S   e r r o r  
    
     r u n t i m e   e r r o r       R u n t i m e   E r r o r ! 
 
 P r o g r a m :     < p r o g r a m   n a m e   u n k n o w n >     . . .   
 
         M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y         atan2        �x��UUU��U��������xx��&�   �   �    �   (�   8�   @�   H�   P�	   X�
   `�   h�   p�   x�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ȸ   и   ظ   �   �   �   ��    �    �!   �"   �#    �$   (�%   0�&   8�'   @�)   H�*   P�+   X�,   `�-   h�/   p�6   x�7   ��8   ��9   ��>   ��?   ��@   ��A   ��C   ��D   ��F   ȹG   йI   عJ   �K   �N   �O   ��P    �V   �W   �Z   �e    �   (�  ,�  8�  D�  P�  \�  h�  t�  ��	  ��  ��  ��  ��  ��  Ⱥ  Ժ  �  �  ��  �  �  �  (�  4�  @�  L�  X�  d�  p�  |�   ��!  ��"  ��#  ��$  ��%  Ļ&  л'  ܻ)  �*  ��+   �,  �-  $�/  0�2  <�4  H�5  T�6  `�7  l�8  x�9  ��:  ��;  ��>  ��?  ��@  ��A  ̼C  ؼD  �E  ��F  �G  �I   �J  ,�K  8�L  D�N  P�O  \�P  h�R  t�V  ��W  ��Z  ��e  ��k  ��l  ̽�  ؽ  �  �  ��	  �
  �   �  ,�  8�  D�  P�  \�  t�,  ��;  ��>  ��C  ��k  Ⱦ  ؾ  �  �	  ��
  �  �   �;  8�k  D�  T�  `�  l�	  x�
  ��  ��  ��;  ��  ��  Ŀ  п	  ܿ
  �  ��   �;  �  (�	  4�
  @�  L�  X�;  p�  ��	  ��
  ��  ��;  ��   ��	   ��
   ��;   ��$   �	$  �
$  �;$  $�(  4�	(  @�
(  L�,  X�	,  d�
,  p�0  |�	0  ��
0  ��4  ��	4  ��
4  ��8  ��
8  ��<  ��
<  ��@  ��
@   �
D  �
H  �
L  $�
P  0�|  <�|  L�(�B   x�,   T�q   �    `��   l��   x��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��C   ���   ��   ��   `�)    ��   8�k    �!   P�c   �   \�D   h�}   t��    �   ��E   8�   ��G   ���   @�   ��H   H�   ���   ���   ��I   ���   ���    �A   ���   P�   �J   X�   ��    ��   ,��   8��   D��   P��   \��   h��   t��   ���   ��K   ���   ���   `�	   ���   ���   ���   ���   ���   ���   ���   ��   ��   ��   (��   4��   @��   L��   X��   d��   p��   |��   ���   0�#   ��e   h�*   ��l   H�&   ��h   h�
   ��L   ��.   ��s   p�   ���   ���   ���   ��M    ��   ��   �>   ��   й7   $�   x�   0�N   ��/   <�t   ظ   H��   T�Z   ��   `�O   X�(   l�j   �   x�a   ��   ��P   ��   ���   ��Q   ��   ��R   ��-   ��r   ��1   ��x   �:   ���   ��   �?   ���   ��S   ��2   ��y   @�%    �g   8�$   �f   ��   p�+   $�m   0��    �=   <��   �;   H��   ��0   T��   `�w   l�u   x�U   ��   ���   ��T   ���   ��   ���   ȹ6   ��~   ��   ��V   ��   ��W   ���   ���   ���   ��   ȸ   �X   и    �Y   ��<   ,��   8��   D�v   P��   �   \�[   (�"   h�d   t��   ���   ���   ���   ���   ���   �   ��\   L��   ���   ���   ��   (��   �   @��   L�]   ��3   X�z   �@   d��   ع8   t��   �9   ���   ��   ��^   ��n    �   ��_   ��5   ��|   �    ��b   �   ��`   ��4   ���   ��{   P�'   �i   �o   �   ,��   <��   H��   T��   `��   l�F   x�p   a r     b g     c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     u k     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k   s y r   d i v       a r - S A   b g - B G   c a - E S   z h - T W   c s - C Z   d a - D K   d e - D E   e l - G R   e n - U S   f i - F I   f r - F R   h e - I L   h u - H U   i s - I S   i t - I T   j a - J P   k o - K R   n l - N L   n b - N O   p l - P L   p t - B R   r o - R O   r u - R U   h r - H R   s k - S K   s q - A L   s v - S E   t h - T H   t r - T R   u r - P K   i d - I D   u k - U A   b e - B Y   s l - S I   e t - E E   l v - L V   l t - L T   f a - I R   v i - V N   h y - A M   a z - A Z - L a t n     e u - E S   m k - M K   t n - Z A   x h - Z A   z u - Z A   a f - Z A   k a - G E   f o - F O   h i - I N   m t - M T   s e - N O   m s - M Y   k k - K Z   k y - K G   s w - K E   u z - U Z - L a t n     t t - R U   b n - I N   p a - I N   g u - I N   t a - I N   t e - I N   k n - I N   m l - I N   m r - I N   s a - I N   m n - M N   c y - G B   g l - E S   k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A   m i - N Z   a r - I Q   z h - C N   d e - C H   e n - G B   e s - M X   f r - B E   i t - C H   n l - B E   n n - N O   p t - P T   s r - S P - L a t n     s v - F I   a z - A Z - C y r l     s e - S E   m s - B N   u z - U Z - C y r l     q u z - E C     a r - E G   z h - H K   d e - A T   e n - A U   e s - E S   f r - C A   s r - S P - C y r l     s e - F I   q u z - P E     a r - L Y   z h - S G   d e - L U   e n - C A   e s - G T   f r - C H   h r - B A   s m j - N O     a r - D Z   z h - M O   d e - L I   e n - N Z   e s - C R   f r - L U   b s - B A - L a t n     s m j - S E     a r - M A   e n - I E   e s - P A   f r - M C   s r - B A - L a t n     s m a - N O     a r - T N   e n - Z A   e s - D O   s r - B A - C y r l     s m a - S E     a r - O M   e n - J M   e s - V E   s m s - F I     a r - Y E   e n - C B   e s - C O   s m n - F I     a r - S Y   e n - B Z   e s - P E   a r - J O   e n - T T   e s - A R   a r - L B   e n - Z W   e s - E C   a r - K W   e n - P H   e s - C L   a r - A E   e s - U Y   a r - B H   e s - P Y   a r - Q A   e s - B O   e s - S V   e s - H N   e s - N I   e s - P R   z h - C H T     s r     a f - z a   a r - a e   a r - b h   a r - d z   a r - e g   a r - i q   a r - j o   a r - k w   a r - l b   a r - l y   a r - m a   a r - o m   a r - q a   a r - s a   a r - s y   a r - t n   a r - y e   a z - a z - c y r l     a z - a z - l a t n     b e - b y   b g - b g   b n - i n   b s - b a - l a t n     c a - e s   c s - c z   c y - g b   d a - d k   d e - a t   d e - c h   d e - d e   d e - l i   d e - l u   d i v - m v     e l - g r   e n - a u   e n - b z   e n - c a   e n - c b   e n - g b   e n - i e   e n - j m   e n - n z   e n - p h   e n - t t   e n - u s   e n - z a   e n - z w   e s - a r   e s - b o   e s - c l   e s - c o   e s - c r   e s - d o   e s - e c   e s - e s   e s - g t   e s - h n   e s - m x   e s - n i   e s - p a   e s - p e   e s - p r   e s - p y   e s - s v   e s - u y   e s - v e   e t - e e   e u - e s   f a - i r   f i - f i   f o - f o   f r - b e   f r - c a   f r - c h   f r - f r   f r - l u   f r - m c   g l - e s   g u - i n   h e - i l   h i - i n   h r - b a   h r - h r   h u - h u   h y - a m   i d - i d   i s - i s   i t - c h   i t - i t   j a - j p   k a - g e   k k - k z   k n - i n   k o k - i n     k o - k r   k y - k g   l t - l t   l v - l v   m i - n z   m k - m k   m l - i n   m n - m n   m r - i n   m s - b n   m s - m y   m t - m t   n b - n o   n l - b e   n l - n l   n n - n o   n s - z a   p a - i n   p l - p l   p t - b r   p t - p t   q u z - b o     q u z - e c     q u z - p e     r o - r o   r u - r u   s a - i n   s e - f i   s e - n o   s e - s e   s k - s k   s l - s i   s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l   s r - b a - c y r l     s r - b a - l a t n     s r - s p - c y r l     s r - s p - l a t n     s v - f i   s v - s e   s w - k e   s y r - s y     t a - i n   t e - i n   t h - t h   t n - z a   t r - t r   t t - r u   u k - u a   u r - p k   u z - u z - c y r l     u z - u z - l a t n     v i - v n   x h - z a   z h - c h s     z h - c h t     z h - c n   z h - h k   z h - m o   z h - s g   z h - t w   z u - z a       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       ���P�Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy HH:mm:ss    S u n   M o n   T u e   W e d   T h u   F r i   S a t   S u n d a y     M o n d a y     T u e s d a y   W e d n e s d a y   T h u r s d a y     F r i d a y     S a t u r d a y     J a n   F e b   M a r   A p r   M a y   J u n   J u l   A u g   S e p   O c t   N o v   D e c   J a n u a r y   F e b r u a r y     M a r c h   A p r i l   J u n e     J u l y     A u g u s t     S e p t e m b e r   O c t o b e r   N o v e m b e r     D e c e m b e r     A M     P M     M M / d d / y y     d d d d ,   M M M M   d d ,   y y y y   H H : m m : s s                       8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7      �?5�h!���>@�������             ��      �@      �                          �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC                                            �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               �       �      ��      ������    ����    ��      ��            8C      8C      0<      0<��+eGW@��+eGW@  ��B.�?  ��B.�?:;����=:;����=�ѱt�?Z�fUUU�?���&WU�?{������?                Mu�{�<`�w>�,  �g5RҌ<t�ӰY  a��aN�`<țuE�  l{�]���<��lX�  ќ/p=�><���2��  ؼcnQ�<P[� {8�&TŤ<�-���B �?RbSQ�<zQ}<�r �S?���<u�o�[� _/:>��<��h1�� �æDAo�<֌b�; �������<8bunz8 ���+G�<�|�eEk 1�	m���<����� �
r�7�<䦅� ���MuM�<�1
� J��]9ݏ<�d�< )}̌/�<ʩ:7�q �^�s)ҧ<���4ۧ mL*�H��<"4L�� ��%F��<).�!
 ��`�cC<-�a`N y����n<�<���� ��z�ΐv<'*6�ڿ 	*(�̃�<�,�v�� ���	�<�O�V+4 ���5�<�'�6Go 	T��c�<)TH�� 5�d+�2�<H!�o� 
���<�U:�~$ �s ��<$"U�8b qU�M��<�;f�� �GΆ�+�<.e<�� �o � �<s_��u ���"a�<�gBV�_ ��F�D�<��s� Ul֫��e<bN�6�� �g�����<�L��% ���<�D��h ����/��<۠*B� D_�Y��{<6w��� <(��`�<��Ͱ77	 �b� ��<ONޟ�}	 'Α+��q<�𣂑�	 �.�X4m�<d�]{f
 ����|'�<\%>�U
 �Zsn�i�<��yUk�
 �3˒w�<��Z���
 �-�f$�<�O��3 ���.�<F^��v ��_
��t<��K�� ��0�ns<�R�ݛ �Y	я��<K�W.�g h�l,kg<i��� � ���6	p�<{�J- �=���t<����X ����PZ�<�2�� ��Js��<^�{3�� ӈ:`�t<�?��.P &I	�'o�<ِ����  �A�Î<'Za�� ��1�d�<@En[vP �͑M;�w<ؐ����       �?       �9��B.�@  ׽2b      �        �������         0<  0<�dW�dW       ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          q7�����8            �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �sinh    cosh    tanh    atan2   fabs    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter  �9:::(:4:@:P:\:d:l:x:�:x��:�:�:�:�:�:�:�:�:�:�:�:�:�:���:�:�:�:���:�:�:�:�:�:t� ;;;;;;;; ;$;(;,;0;4;8;D;P;X;d;|;�;�;�;�;�;<<<`<|<�<�<�<=== =0=T=\=h=x=�=�=�=>,>X>t>�>�>�>?x�0?D?`?t?�?__based(    __cdecl __pascal    __stdcall   __thiscall  __fastcall  __vectorcall    __clrcall   __eabi  __ptr64 __restrict  __unaligned restrict(    new     delete =   >>  <<  !   ==  !=  []  operator    ->  *   ++  --  +   &   ->* /   <   <=  >   >=  ,   ()  ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall' `typeof'    `local static guard'    `string'    `vbase destructor'  `vector deleting destructor'    `default constructor closure'   `scalar deleting destructor'    `vector constructor iterator'   `vector destructor iterator'    `vector vbase constructor iterator' `virtual displacement map'  `eh vector constructor iterator'    `eh vector destructor iterator' `eh vector vbase constructor iterator'  `copy constructor closure'  `udt returning' `EH `RTTI   `local vftable' `local vftable constructor closure'  new[]   delete[]   `omni callsig'  `placement delete closure'  `placement delete[] closure'    `managed vector constructor iterator'   `managed vector destructor iterator'    `eh vector copy constructor iterator'   `eh vector vbase copy constructor iterator' `dynamic initializer for '  `dynamic atexit destructor for '    `vector copy constructor iterator'  `vector vbase copy constructor iterator'    `managed vector copy constructor iterator'  `local static thread guard'  Type Descriptor'    Base Class Descriptor at (  Base Class Array'   Class Hierarchy Descriptor'     Complete Object Locator'   U S E R 3 2 . D L L     MessageBoxW GetActiveWindow GetLastActivePopup  GetUserObjectInformationW   GetProcessWindowStation           8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �        ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               ( ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                                                            �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#SNAN  1#IND   1#INF   1#QNAN  C O N O U T $   A      H                                                           �`�   RSDS�I>�@?DB�����|�   E:\repos\cmNodes\src\obj\cmnodes_r13_Win32_Release.pdb      �   �                      �j�j�j    X�       ����    @   |jp�        ����    @   �j           �j�j               �jk�j    ��       ����    @   �j            ��4k           DkPk�j    ��       ����    @   4k           |k�k�j�j    ��       ����    @   lk           �k�k�j�j    ܲ       ����    @   �k��       ����    @    l           l�k lXl    �       ����    @   <l           Ll lXl    ,�        ����    @   tl           �lXl                D��l           �l�l�l    D�       ����    @   �l`�        ����    @   �l           m�l                |� m           0mDm�k lXl    |�       ����    @    m            ��tm           �m�mk�j    ��       ����    @   tm            ���m           �m�mn�j�j    ��       ����    @   �mȳ       ����    @    n           0nn�j�j                �Tn           dnxnn�j�j    �       ����    @   Tn            ��n           �n�n�j�j    �       ����    @   �n            (��n           oo�k�j�j    (�       ����    @   �n            D�Lo           \opo�o�j�j    D�       ����    @   Lo`�       ����    @   �o           �o�o�j�j                |��o           �o p�o�j�j    |�       ����    @   �o            ��0p           @pTp�o�j�j    ��       ����    @   0p            ���p           �p�p�o�j�j    ��       ����    @   �p            Դ�p           �p�p�o�j�j    Դ       ����    @   �p            �,q           <qPq�o�j�j    �       ����    @   ,q            ��q           �q�q�o�j�j    �       ����    @   �q            (��q           �q�q�o�j�j    (�       ����    @   �q            D�(r           8rLr�o�j�j    D�       ����    @   (r            `�|r           �r�r�o�j�j    `�       ����    @   |r            |��r           �r�r�o�j�j    |�       ����    @   �r            ��$s           4sHs�o�j�j    ��       ����    @   $s            ��xs           �s�s�o�j�j    ��       ����    @   xs            Ե�s           �s�s�o�j�j    Ե       ����    @   �s            �� t           0tDt�o�j�j    ��       ����    @    t            �tt           �t�t�o�j�j    �       ����    @   tt            0��t           �t�t�o�j�j    0�       ����    @   �t            L�u           ,u@u�o�j�j    L�       ����    @   u            h�pu           �u�u�o�j�j    h�       ����    @   pu            ���u           �u�u�o�j�j    ��       ����    @   �u            ��v           (v<v�o�j�j    ��       ����    @   v            ��lv           |v�v�o�j�j    ��       ����    @   lv            ܶ�v           �v�v�o�j�j    ܶ       ����    @   �v            ��w           $w8w�o�j�j    ��       ����    @   w            �hw           xw�w�o�j�j    �       ����    @   hw            8��w           �w�w�o�j�j    8�       ����    @   �w            X�x            x4x�o�j�j    X�       ����    @   x            t�dx           tx�x�o�j�j    t�       ����    @   dx            ���x           �x�x�o�j�j    ��       ����    @   �x            ��y           y0y�o�j�j    ��       ����    @   y            ̷`y           py�y�o�j�j    ̷       ����    @   `y            ��y           �y�y�o�j�j    �       ����    @   �y            �z           z,z�o�j�j    �       ����    @   z             �\z           lz�z�o�j�j     �       ����    @   \z            @��z           �z�z�o�j�j    @�       ����    @   �z            `�{           {({�o�j�j    `�       ����    @   {            ��X{           h{|{�o�j�j    ��       ����    @   X{            ���{           �{�{Pk�j    ��       ����    @   �{            ���{           ||Pk�j    ��       ����    @   �{            �L|           \|l|Pk�j    �       ����    @   L|             ��|           �|�|Pk�j     �       ����    @   �|             ��|           �|}Pk�j     �       ����    @   �|            D�<}           L}\}Pk�j    D�       ����    @   <}            h��}           �}�}Pk�j    h�       ����    @   �}            ���}           �}�}Pk�j    ��       ����    @   �}            ��,~           <~L~Pk�j    ��       ����    @   ,~            Թ|~           �~�~Pk�j    Թ       ����    @   |~            ���~           �~�~Pk�j    ��       ����    @   �~            �           ,<Pk�j    �       ����    @               <�l           |�Pk�j    <�       ����    @   l            \��           ��Pk�j    \�       ����    @   �            |��           �,�Pk�j    |�       ����    @   �            ��\�           l�|�Pk�j    ��       ����    @   \�            ����           ��̀Pk�j    ��       ����    @   ��            ���           ��Pk�j    �       ����    @   ��            �L�           \�l�Pk�j    �       ����    @   L�            @���           ����Pk�j    @�       ����    @   ��            h��           ���Pk�j    h�       ����    @   �            ��<�           L�\�Pk�j    ��       ����    @   <�            Ļ��           ����Pk�j    Ļ       ����    @   ��            �܂           ���Pk�j    �       ����    @   ܂            �,�           <�L�Pk�j    �       ����    @   ,�            @�|�           ����Pk�j    @�       ����    @   |�            h�̃           ܃�Pk�j    h�       ����    @   ̃            ���           ,�<�Pk�j    ��       ����    @   �            ��l�           |���Pk�j    ��       ����    @   l�            ���           ̄܄Pk�j    �       ����    @   ��            ��           �,�Pk�j    �       ����    @   �            <�\�           l�|�Pk�j    <�       ����    @   \�            l���           ��̅Pk�j    l�       ����    @   ��            ����           ��Pk�j    ��       ����    @   ��            ĽL�           \�l�Pk�j    Ľ       ����    @   L�            ���           ����Pk�j    �       ����    @   ��            ��           ���Pk�j    �       ����    @   �            H�<�           L�\�Pk�j    H�       ����    @   <�            t���           ����Pk�j    t�       ����    @   ��            ��܇           ���Pk�j    ��       ����    @   ܇            Ⱦ,�           <�L�Pk�j    Ⱦ       ����    @   ,�            ��|�           ����Pk�j    ��       ����    @   |�             �̈           ܈�Pk�j     �       ����    @   ̈            L��           ,�<�Pk�j    L�       ����    @   �            x�l�           |���Pk�j    x�       ����    @   l�            ����           ̉܉Pk�j    ��       ����    @   ��            Կ�           �,�Pk�j    Կ       ����    @   �            �\�           l�|�Pk�j    �       ����    @   \�            ,���           ��̊Pk�j    ,�       ����    @   ��            X���           ��Pk�j    X�       ����    @   ��            ��L�           \�l�Pk�j    ��       ����    @   L�            ����           ����Pk�j    ��       ����    @   ��            ���           ���Pk�j    ��       ����    @   �            �<�           L�\�Pk�j    �       ����    @   <�            0���           ����Pk�j    0�       ����    @   ��           ،�Pk�j    X�       ����    @   Ȍ            ���           (�<��Pk�j    ��       ����    @   �            ��l�           |����Pk�j    ��       ����    @   l�            ����           Ѝ��Pk�j    ��       ����    @   ��            ��           $�8��Pk�j    �       ����    @   �            4�h�           x����Pk�j    4�       ����    @   h�            `���           ̎���Pk�j    `�       ����    @   ��            ���            �4��Pk�j    ��       ����    @   �            ��d�           t����Pk�j    ��       ����    @   d�            ����           ȏ܏�Pk�j    ��       ����    @   ��            ��           �0��Pk�j    �       ����    @   �            <�`�           p�|��l    <�       ����    @   `�            `���           ��ȐXl    `�       ����    @   ��            ����           ��Pk�j    ��       ����    @   ��            ��H�           X�d�Xl    ��       ����    @   H�            ����           ����Pk�j    ��       ����    @   ��            ���           �� ��    ��       ����    @   ��        ����    @   8�           H��                ,�d�           t����k�j�j    ,�       ����    @   d�            `��o            p��j            �8�            �<l            ,�tl            `��l            H�0�           @�L�Xl    H�       ����    @   0�            �� l            d���           ����    d�        ����    @   ��           ԓܓ    |�        ����    @   ē            ���           �(�ܓ    ��       ����    @   �            ��X�           h�p�    ��        ����    @   X�            ����           ����p�    ��       ����    @   ��            ȳ n            �� �           ��    ��        ����    @    �            �H�           X�`�    �        ����    @   H�            0���           ����    0�        ����    @   ��            P�ؕ           ���ܓ    P�       ����    @   ؕ            t�$�           4�<�    t�        ����    @   $�        �  T ��                     ����    ����    ����    �    ����    ����    ��������    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    W�����    c�����    ����    ����    ������    ������    ����    ����    H�    ����    |���    ����    %�    ����    ����    ����    �    ����    ����    ����    M    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    @!    ����    ����    ����    �"    ����    ����    �����P�P    ����    ����    ����    *S    ����    ����    �����cd    ����    ����    �����d�d    ����    ����    ����    �r    ����    ����    ����    at        +t����    ����    ����    �t    ����    ����    ����    т    ����    ����    ����    Q�    ����    ����    ����    !�    ����    ����    ����    �                ߃DT    �          � � � J �   cmnodes_r13.cdl c4d_main  4�         ��  �                     ,� <� L� ^� t� �� �� �� �� ̛ ܛ �  � � (� >� P� `� n� �� �� �� Ȝ ޜ �� � ,� H� f� �� �� �� �� ʝ ؝ � � � � &� 2� B� Z� r� �� �� �� �� Ğ О ܞ � �� � � 0� @� P� b� v� ��     !EncodePointer � DecodePointer �GetCommandLineA GetCurrentThreadId  PGetLastError  3HeapFree  /HeapAlloc mIsProcessorFeaturePresent gIsDebuggerPresent 
SetLastError  QExitProcess fGetModuleHandleExW  �GetProcAddress  �MultiByteToWideChar �WideCharToMultiByte �GetProcessHeap  �GetStdHandle  >GetFileType DeleteCriticalSection �GetStartupInfoW bGetModuleFileNameA  -QueryPerformanceCounter 
GetCurrentProcessId �GetSystemTimeAsFileTime 'GetEnvironmentStringsW  �FreeEnvironmentStringsW �UnhandledExceptionFilter  ASetUnhandledExceptionFilter HInitializeCriticalSectionAndSpinCount PSleep 	GetCurrentProcess _TerminateProcess  qTlsAlloc  sTlsGetValue tTlsSetValue rTlsFree gGetModuleHandleW  �WriteFile cGetModuleFileNameW  8HeapSize  �LCMapStringW  %EnterCriticalSection  �LeaveCriticalSection  �GetConsoleCP  �GetConsoleMode  �SetFilePointerEx  rIsValidCodePage �GetACP  �GetOEMCP  �GetCPInfo ?RaiseException  �RtlUnwind �LoadLibraryExW  6HeapReAlloc �OutputDebugStringW   SetStdHandle  �WriteConsoleW �GetStringTypeW  �FlushFileBuffers  � CreateFileW  CloseHandle KERNEL32.dll                                                                                                                 N�@���Du�  s�     ����                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                acos            atan            cos                   �?pow     sin             sqrt    ?  ?  cccccccccc����    �����
                                                          ����            asin            log     ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                            0��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��               C   ������ ������ �(�4�@�H�T�X�\�`�d�h�l�p�t�x�|�����������d��������������������� ��        �(�0�8�@�H�P�X�h�x�������������������������$�,�4�D�X�d���p�|������������������0�����                                   T�            T�            T�            T�            T�                          خ        b�fhX�                        �����&     �   �   ��   ��    8   8!   8   �   �   $�   8   P�   D�   H�    L�   ,�   4�    8   <�   (8   08   88   @8   H8"   P8#   T8$   X8%   \8&   d8      �      ���������              �       �D        � 0                                                                                                                                                                                                                                                                                           خ.   Ԯ������������������(���������������.   bd             �            d   ���5      @   �  �   ����             ����         �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                  ��`    .?AVNodeData@@  �`    .?AVBaseData@@  �`    .?AVCustomGuiData@@ �`    .?AVCommandData@@   �`    .?AVSceneHookData@@ �`    .?AVShaderData@@    �`    .?AViCustomGui@@    �`    .?AVSubDialog@@ �`    .?AVGeDialog@@  �`    .?AVcmMenuButton@@  �`    .?AVGeUserArea@@    �`    .?AVcmRealDlg@@ �`    .?AVcmRealGui@@ �`    .?AVcmPrefsObject@@ �`    .?AVPrefsDialogObject@@ �`    .?AVcmNodesPrefsObject@@    �`    .?AVcmNodeTree@@    �`    .?AVcmNodeForest@@  �`    .?AVcmNodeOutput@@  �`    .?AVcmNodeBase@@    �`    .?AVcmNodeMaterial@@    �`    .?AVcmNodeTexture@@ �`    .?AVcmNodeColor@@   �`    .?AVcmNodeShuffle@@ �`    .?AVcmNodeCopy@@    �`    .?AVcmNodeBlend@@   �`    .?AVcmNodeMath@@    �`    .?AVcmNodeClamp@@   �`    .?AVcmNodeCurves@@  �`    .?AVcmNodeGrade@@   �`    .?AVcmNodeColorspace@@  �`    .?AVcmNodeFilter@@  �`    .?AVcmNodeColorize@@    �`    .?AVcmNodeInvert@@  �`    .?AVcmNodeTransform@@   �`    .?AVcmNodeDistort@@ �`    .?AVcmNodeEmboss@@  �`    .?AVcmNodeMatrix@@  �`    .?AVcmNodeBlur@@    �`    .?AVcmNodeEdgeDetect@@  �`    .?AVcmNodeDirBlur@@ �`    .?AVcmNodeHighPass@@    �`    .?AVcmNodeInfo@@    �`    .?AVcmNodeSpecular@@    �`    .?AVcmNodeDistance@@    �`    .?AVcmNodeSwitch@@  �`    .?AVcmNodeReflection@@  �`    .?AVcmNodeNoop@@    �`    .?AVcmNodeDiffuse@@ �`    .?AVcmNodeFresnel@@ �`    .?AVcmNodeTiler@@   �`    .?AVcmNodeShadow@@  �`    .?AVcmNodeNormalMap@@   �`    .?AVcmNodeCondition@@   �`    .?AVcmNodeProjector@@   �`    .?AVcmNodeVrayAdvanced@@    �`    .?AVcmNodeCmd_Cut@@ �`    .?AVcmNodeCmd_Copy@@    �`    .?AVcmNodeCmd_Paste@@   �`    .?AVcmNodeCmd_Delete@@  �`    .?AVcmNodeCmd_SelectAll@@   �`    .?AVcmNodeCmd_DeselectAll@@ �`    .?AVcmNodeCmd_Disconnect@@  �`    .?AVcmNodeCmd_FrameSelected@@   �`    .?AVcmNodeCmd_Prefs@@   �`    .?AVcmNodeCmd_AddTree@@ �`    .?AVcmNodeCmd_TreeMenu@@    �`    .?AVcmNodeCmd_NodeMenu@@    �`    .?AVcmNodeCmd_ZoomIn@@  �`    .?AVcmNodeCmd_ZoomOut@@ �`    .?AVcmNodeCmd_Zoom100@@ �`    .?AVcmNodeCmd_ResetView@@   �`    .?AVcmNodeCmd_CalcPreview@@ �`    .?AVcmNodeCreateCmd_NodeSolidColor@@    �`    .?AVcmNodeCreateCmd_NodeTexture@@   �`    .?AVcmNodeCreateCmd_NodeClamp@@ �`    .?AVcmNodeCreateCmd_NodeColorspace@@    �`    .?AVcmNodeCreateCmd_NodeCurves@@    �`    .?AVcmNodeCreateCmd_NodeFilter@@    �`    .?AVcmNodeCreateCmd_NodeGrade@@ �`    .?AVcmNodeCreateCmd_NodeMath@@  �`    .?AVcmNodeCreateCmd_NodeBlend@@ �`    .?AVcmNodeCreateCmd_NodeCopy@@  �`    .?AVcmNodeCreateCmd_NodeShuffle@@   �`    .?AVcmNodeCreateCmd_NodeBlur@@  �`    .?AVcmNodeCreateCmd_NodeDirBlur@@   �`    .?AVcmNodeCreateCmd_NodeDistort@@   �`    .?AVcmNodeCreateCmd_NodeEdgeDetect@@    �`    .?AVcmNodeCreateCmd_NodeEmboss@@    �`    .?AVcmNodeCreateCmd_NodeMatrix@@    �`    .?AVcmNodeCreateCmd_NodeNormalMap@@ �`    .?AVcmNodeCreateCmd_NodeTransform@@ �`    .?AVcmNodeCreateCmd_NodeOutput@@    �`    .?AVcmNodeCreateCmd_NodeMaterial@@  �`    .?AVcmNodeCreateCmd_NodeColorize@@  �`    .?AVcmNodeCreateCmd_NodeInfo@@  �`    .?AVcmNodeCreateCmd_NodeHighPass@@  �`    .?AVcmNodeCreateCmd_NodeSwitch@@    �`    .?AVcmNodeCreateCmd_NodeInvert@@    �`    .?AVcmNodeCreateCmd_NodeSpecular@@  �`    .?AVcmNodeCreateCmd_NodeVrayAdvanced@@  �`    .?AVcmNodeCreateCmd_NodeDistance@@  �`    .?AVcmNodeCreateCmd_NodeReflection@@    �`    .?AVcmNodeCreateCmd_NodeNoop@@  �`    .?AVcmNodeCreateCmd_NodeDiffuse@@   �`    .?AVcmNodeCreateCmd_NodeFresnel@@   �`    .?AVcmNodeCreateCmd_NodeTiler@@ �`    .?AVcmNodeCreateCmd_NodeShadow@@    �`    .?AVcmNodeCreateCmd_NodeCondition@@ �`    .?AVcmNodeCreateCmd_NodeProjector@@ �`    .?AVcmNodeCreateCmd_NodeInput@@ �`    .?AVcmTreeBookmarkCmd_Bookmark@@    �`    .?AVcmTreeBookmarkCmd_Bookmark0@@   �`    .?AVcmTreeBookmarkCmd_Bookmark1@@   �`    .?AVcmTreeBookmarkCmd_Bookmark2@@   �`    .?AVcmTreeBookmarkCmd_Bookmark3@@   �`    .?AVcmTreeBookmarkCmd_Bookmark4@@   �`    .?AVcmTreeBookmarkCmd_Bookmark5@@   �`    .?AVcmTreeBookmarkCmd_Bookmark6@@   �`    .?AVcmTreeBookmarkCmd_Bookmark7@@   �`    .?AVcmTreeBookmarkCmd_Bookmark8@@   �`    .?AVcmTreeBookmarkCmd_Bookmark9@@   �`    .?AVcmNodeEditorUserArea@@  �`    .?AVcmNodeEditorDialog@@    �`    .?AVcmNodeEditorCommand@@   �`    .?AVcmTreeManagerDialog@@   �`    .?AVcmTreeManagerCommand@@  �`    .?AVcmUpdateNodeThread@@    �`    .?AVC4DThread@@ �`    .?AVcmNodeShader@@  �`    .?AVGeModalDialog@@ �`    .?AVNeighbor@@  �`    .?AVGeSortAndSearch@@   �`    .?AVDisjointNgonMesh@@  �`    .?AVGeListView@@    �`    .?AVSimpleListView@@    �`    .?AVGeToolNode2D@@  �`    .?AVGeToolList2D@@  �`    .?AVGeToolDynArray@@    �`    .?AVGeToolDynArraySort@@    �`    .?AVtype_info@@                                                                                                                        0  0$0B0L0T0p0x0�0�0�0�0�0�0�0�0�0�011 141M1^1o1{1�1�1�1�1�1�122$222F2_2|2�2�2�2�2�2�233303I3f3w3�3�3�3�3�3�3�34434P4a4m4{4�4�4�4�4�4�45515B5N5\5t5�5�5�5�5�56%6W6h6�6�6�6�6�6&7c7t7�7�7�7�7�78$888e8�8�8�8�8�8�8
99D9V9`9n9w9�9�9�9�9�9�9�9:-:A:f:p:�:/;c;�=�=�=�=�>�>�>�>?a?i?z?�?�?�?      �   0&0�0�0�01'1�1�1�192J2z2�2�2�2�2;3Q3c3�3�3�3�3�34"4-4;4�56o6�6(7s7�7(8H8�89L9|:�:�:a;�;0<8<�<'=�=�=�>�>7?T?p?�?�?�? 0  �   �0�0�0�0�0�01B1P1[1�1�1�12/2Y2�2�2�2363>3_3�3�3�3�3�4
55D5g5{5�5G6Z6�6�6�6g7�7�7�7�788q9�9�9:�=�=�=>e>�>�>�>+?I?Q?b? @  �   0'090A0L0o0~0�0�0�0�0�0�0�01*1I1`1h1p1�1�12R2�2�2�2�2
3*3>3P3a3y3�3�3�34k4�4�4�4[5~5C6�6�6�6�6�6�6+7g8x8�8�8�8�8�89C9P9e9y9�9�9�9::�:�:�:�:�:;;';e;m;�;�;�;�;�;x<�<�<�<�< =-=B=V=o=�=�=�=�=>	>0>8>K>�?�?�? P  �  0)010U0]0p0�0�0�0�0�0�01
1.1B1J1p1x1�1�1�1�1�1 22#2H2L2P2T2X2\2`2q2�2�2�2�2�2333,3=3R3f3|3�3�3�3�3�34#424C4T4`4�4�4�4�4�4�4�455-5>5J5j5x5�5�5�5�5�5�56$6:6C6`6o6�6�6�6�6�6�6�67"777H7Y7j7{7�7�7�7�7�7�7	88/8@8^8o8{8�8�8�8�8�8�89919T9h9t9�9�9�9�9�9�9::0:A:R:^:x:�:�:�:�:�:�:�:�:;(;A;R;g;{;�;�;�;�;�;<</<@<Q<b<s<<�<�<�<�<�<==&=D=X=d=r=�=�=�=�=�=�=!>.>B>X>b>>�>�>�>�>?/?;?I?Z?f?�?�?�?�?�?   `  L  �0�0�0 11A1[1w1�1�1�1�1�1�1242N2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2N3~3�3�3�3�3454M4`4�4�4�4�4�45%5=5P5s5�5�5�5�5�56-6@6c6{6�6�6�6�6�6707S7k7~7�7�7�7�78+8>8N8c8{8�8�8�8�8�8�89.9F9Y9�9�9�9�9�9�9:(:>:N:c:{:�:�:�:�:�:�:;;3;K;`;v;�;�;�;�;�;�;<<�<=;=[=�=�=�=�=�=�=�=�=�=>6>G>S>a>u>�>�>�>�>�>?A?G?r?~?�?�?�?�?   p  (  !080E0O0�0�0�0�0�0�0111:1V1g1p1�1�1�1�1�1�1�12 2)2:2F2T2e2q2�2�2�2�2�2�233)3:3C3_3p3y3�3�3�3�3�3�3�34434G4X4k4t4�4�4�4�4�4�4�4�4	5.5B5S5f5o5�5�5�5�5�5�5�5�56(696E6S6d6p6�6�6�6�6�6�677(797B7^7o7x7�7�7�7+:K:�:�:;S;m;�;�;�;�;�;�;�; <#</<C<d<y<�<�<4=[=o=�=�=�=�=$>_>�>�>?,?D?�?�?   �  `  T0�0�0�0d1x1�1�1�1�1�1�1�1	22+2@2T2v2�2�2�2�2�2�233C3T3e3�3�3�3�3�3�3'484I4Z4u4�4�4�4�4�4	5.5?5^5s5�5�5�5�5�56662686]6g6{6�6�6�6�6�6�6�6�6�67%7T7i7u7�7�7�7�7�7�78*8;8O8e8v8�8�8�8�8�8�89 9=9Y9j9v9�9�9�9�9�9::1:O:`:y:�:�:�:�:�:	;';8;Q;o;�;�;�;�;�;�;<)<G<X<q<�<�<�<�<�<==0=I=g=x=�=�=�=�=�=>!>?>P>i>�>�>�>�>�>�>?(?A?_?p?�?�?�?�?�?   �     0070H0a00�0�0�0�0�01 191W1h1�1�1�1�1�1�12/2@2Y2w2�2�2�2�2�23313O3`3y3�3�3�3�3�344+4k4|4�4�4�4�4�4�4�4;5L5]5w5�5�5�5�5�5�5�56626L6b6~6�6�6�6�6�6�67)7:7x7�7�7�78%8b8n8�8�89*9]9�9�9�9�9�9:";*;8;T;b;n;|;�;�;�;�;�;�;<,<{<�<�<�<=-=A=|=�=�=�=�=�=�=�=�=�=>*?6?U?k?   �  �   �2�2�2�2�3�3�3484h4�4�485h5�5�5�5(6X6�6�6H7x7�7�7�7 888h8�8�8�8(9X9�9�9�9:H:x:�:�:;8;k;t;�;�;<H<�<�<(=\=j=v=�=�=> >1>=>[>p>�>�>??+?3?R?\?z?�?�?�?�?�? �  8  0$0B0I0i0�0�0�0�0�0	121<1\1�1�1�1�1�12#2B2L2j2v2�2�2�2�2�2"3,3K3S3r3|3�3�3�3�3�3�344:4F4b4l4�4�4�4�455+535R5\5}5�5�5�5�56"6)6I6X6�6�6�6�6�6�67	7(707Q7[7�7�7�7�7�7�7�78868Q8[8�8�8�8�8�8�8929<9[9c9�9�9�9�9�9
::R:\:y:�:�:�:�:�:�:;;<;R;];r;y;�;�;�;�;�;�;<2<9<V<v<}<�<�<= =,=H=�=�=>$>�>�>�>�> �  �   i1z1�1�1O2`2l2�2�2�2�2�2�23303A3R3^33�3�3�3�3�3�34"434D4P4q4�4�4�4�4�4�4�45 515=5^5y5�5�5�5�5�5�56�6T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7 88888888 8$8(8>8�8�8�8�8�8�8�8�8�8�8�8�8�8�89?9a9�9�9: :�;�;%=)>w>�? �  �   '0�0�0�0�0121S1h1�1222`2�2�2�2-5�5�6�6�6�7)8M8�8�8�8�8�8�809L9h9�9 : :�:�:�:�:w;�;<;<J<p<�<�<D=S=y=�=#>+>9>L>�>�>�>�>�>?3?D?�?   �  �    00040�0�0�0�0�0�0 1111181I1U1c1�1�1�1�1�1�1�1	232D2P2^2e3�3�3�3�3/4@4L4Z4v4�4�4�4�4�4�45+5R5i5�5�5�5�56+6W6k6�6787}7�7�7�7�7�7�78(848B8S8�8�8�8999a9{9�9�9�9*:J:k:�:�:�:;; ;4;b;�;�;�;�;�;�;%<H<�<�<�<=5=O=�=�=�=�=>8>I>x>�?�?   �  ,  00�0�0�0�0�011'1k1�1�1222h2y2�2�2�2�2#3�3�3�3�3�3�3�3�3�3�3X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56&6/6N6_6p6|6�6G7X7d7�7�7�7�78O8`8l8�8999=9N9_9k9�9:M:h:q:�:�:�:�:�:;;!;/;Y;j;v;�;�;�;�;�;A<a<�<�<�<-=M=�=�=�=>!>=>^>�>�>�>4?C?a?�?�?     h  0_0p0�0�0%1g1x1�1�1�1J2j2�23W3i3�3�3�3�3�3�34C4T4`4n4�4�4�4�4�4�4X5i5u5�5�5#646@6N6b6�6�6�6�67X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;<�<�<�<�<_=p=|=�=�=�>�>�>�>?"?.?<?�?�?  `   0+0~12�2�23(3�34Z4c4s4�4�455E5X5�5�516�6�7�7�8�8�; <Z<g<�<=�=�=:>K>W>p>�>�>??F?   �   ,0L0m0�0�0�0�0�011$2�2�2373u3�3�3�344N4_4�4�4�4�45F6R6�6�6�6�6�6�6}7�7�7�7�7s8�8�9�9
::?:`:s:�:�:�:;;5;�;<4<F<v<�<�<=6=R=h=�=>b>�>H?^?�?�?   0 �   000!0.0[0~0�0�0 111#1�1�1%282�2�2�2�2�23Q3d3�3�3r4�4�455�5�56L67$7Y7a7�7�7]859I9�9�9.:�:�:*;?;�;q<�<�<�<!=.=�>�>   @ X   a0�0�1�12e2�23\3�:�:;z;�;�;�;�;�;<#<4<E<V<�<�<�<�<==V=g=x=�=�=>7>P>c>??G? P �   90q0�0�01!1&171C1Q1c1�1�1�1�1�1�1�1�12242E2Q2_2r2�2�2�2�2�23,3w4�4�4�4�4O5i5�5�576Q6�6�6797�7�78!8{8�8�8	9c9}9�9�9K:e:�:�:3;M;�;�;<h<�<�<�<=u=�=>%>n>�>�>%?n?�?�?�? ` �   0,0J0}0�0�01111%1n1�1�1�1�2�2�2�233/3B3a3j3y3�3444�4�45%545I5i5�5�5�5�5	6O6e6t6�6�6�677)7I7�7�7�7�7�7/8E8T8i8�8�8�8d9�9�9�9 :Q:�:N;U;Z;k;�;�;�;*<;<�<�<�<�<�<=1=N=k=�=�=�=�=>>>>>>> >$>(>,>�>�>�>+?X?�?�?�?   p d  090f0�0�0�01G1t1�1�1�1(2U2�2�2�2	363c3�3�3�34D4q4�4�4�4%5R55�5�5636`6�6�6�67A7n7�7�7�7"8O8|8�8�8909]9�9�9�9:>:k:�:�:�:7;T;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<=,=>=G=�=�=�=�=�=>%>,>>>D>o>~>�>�>�>�>&?8???Q?X?j?p?�?�?�?�?�? � �  	0 070N0e0|0�0�0�0�0�0�0�0�0�0�0�0�01(1/1A1H1Z1`1�1�1�1�1�122"262H2Y2j2|2�2�2�2$353A3O3e3y3�3�3�3�3�3�3�3M4\4e4�4�4�4�4�4�45'5>5U5l5�5�5�5�5�5�56$6;6R6i6�6�6�6�6�6�6
7!787O7f7}7�7�7�7�7�78858L8c8z8�8�8�8�8�89929I9`9w9�9�9�9�9�9::/:F:]:t:�:�:�:�:�:�:;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<g<�<�<�<1=h=�=�=�=7>�>�>�>�> ???-?j?�?�?�? � �   00�0�01!1H1a1�1�1�112i2�2�2�233*3@3Y3o3�3�3�3�3�3�3 44&4:4S4d4y4�4�4�4�4�4�4�4!5D5t5�5�5A6�6�677�7�7�7�7�78�8�8�8�89;9:!:J:e:�:8;�;�;�;�;�;�;<<!<<<n<}<�<�<�<�<�<�<�<=Q=`={=�=�=�=�=�=�=,>=>t>�>�>�>�>�><?f?�?�?�?�?   � H  0#0/0=0X0�0�0�0�0161T1�1�1�1�1�12!2Q2�2�2�2�2�2.3=3G3a3l3�3�3�3�3�3�3404F4Q4j4�4�4�4�45,5K5V5o5z5�5�5�5�5�56616^6m6w6�6�6�6�677<7[7z7�7�7�7�7�78'828d8}8�8�8�8�89999O9e9�9�9�9�9�9�9�9:.:9:R:]:v:�:�:�:�:�:�:;';a;p;�;�;�;�;�;�;	<<&<4<O<�<�<�<�<�<�<='===S=i==�=�=�=�=> >1>=>K>f>�>�>�>�>�>?/?^?m?w?�?�?�?�? � @   0020H0g0�0�0�0�0�0�0�0
1$1I1�1�1�1�1�1�1282`2~2�2�2�2�23>3M3i33�3�3�3�3�34$4:4P4�4�4�4�4�4�4�4.5=5Y5o5�5�5�5�5�5�56686C6~6�6�6�6�6�677-7C7Y7o7�7�7�7�7�7�7	8858K8a8w8�8�8�8�8�8�89'9=9S9i99�9�9�9�9�9::/:E:[:q:�:�:�:�:�:�:;!;7;M;c;y;�;�;�;�;�;�;<)<?<U<k<�<�<�<�<�<�<==1=G=]=s=�=�=�=�=�=�=>#>�?   � �   �0X1\1`1d1h1l1p1t1�1�1�1252S2�2�23M3�3D4�45�56t6�6�6D7^7r7�7�7�748F8�8�8�89H9i9z9�9�9�9�9:::-:T:x:�:�:�:�:�:�:(;X;i;u;�;�;�;�;<<!</<�<�<�<�=�=�=�=9>W>�>�>�>�> � �   
0A0�0�0�0�0�0�0A1|1�1�1�1�12F2Q2�23H3�3�3�3�3�3�3*4q4�4�4�4�45D5h5�5�5�5�5�5t6�6{7�7�7�7�7�788(8D8c8m8�8�8�8�8�899/9K9^9w9�9�9�9�9�;�;�<D>d>h>l>p>t>x>|>�>�>�>�>?�?�?   � l   0?0q1�1K2\2h2v2�2�2�2�2�233'3[3l3x3�3�34�5�5�5�6�6�6�6788:':�=�=�=>G>i>z>�>�>�>�>?? ?b?�? � �  00[0�0�0�0�0�0�0�0111@1N1�1�1�2�2�2�2�2�2 3/3U3w3�3�3�344&4?4X4i4�4�4�4�4�4�45505D5�5�5�5�5�5�5�5�5 66666t6x6|6�6�6�6�6�6�6�6�6�6�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9$:8:J:Q:n:w:�:�:�:�:�:�:�:;;1;B;Z;k;�;�;�;�;�;�;4<H<Z<d<�<�<�<�<�<�<�<�<==+=D=U=m=~=�=�=�=�= >>D>X>j>q>�>�>�>�>�>�>�>??$?8?Q?b?z?�?�?�?�?�?   �  00T0h0z0�0�0�0�0�0�0�0�01141H1a1r1�1�1�1�1�122.2d2x2�2�2�2�2�2�2�2�2�2"3/3D3X3q3�3�3�3�3�344-4>4t4�4�4�4�4�4�4�4�45525?5T5h5�5�5�5�5�5�56,6=6N6�6�6�6�6�6�6�6�6777B7O7d7x7�7�7�7�7�78+8<8M8^8�8�8�8�8�8�8�899#9/9R9_9t9�9�9�9�9�9::;:L:]:n:�:�:�:�:�:�:;;%;6;B;e;r;�;�;�;�;�;�;<2<N<_<p<�<�<�<�<�<�<==$=2=C=O=r==�=�=�=�=�=�=+>?>[>l>}>�>�>�>�>�>??(?4?B?S?_?�?�?�?�?�?�?�?    �  0;0O0k0|0�0�0�0�0�01!1*1;1G1U1f1r1�1�1�1�1�1�122N2b2~2�2�2�2�2�2
33.373H3T3b3s33�3�3�3�3�344+4[4o4�4�4�4�4�455$5A5J5[5g5u5�5�5�5�5�5�566-6>6n6�6�6�6�6�677*747Q7Z7k7w7�7�7�7�7�7�7�78%8=8N8~8�8�8�8�8�89(9:9D9a9j9{9�9�9�9�9�9�9�9:$:5:M:^:�:�:�:�:�:�:$;8;J;T;q;z;�;�;�;�;�;�;�;<<4<E<]<n<�<�<�<�<�<=3=G=Y=c=�=�=�=�=�=�=�=�=�=�=
>>3>G>`>q>�>�>�>�>	??+?<?s?�?�?�?�?�?�?�?�?   �  00000<0J0[0s0�0�0�0�0�0'181I1Z1k1|1�1�1�1�1 2	22&242E2Q2_2p2|2�2�2�2�2�2�233g3x3�3�3�3�3�344#4@4I4Z4f4t4�4�4�4�4�4�4�4�45 515F5Z5�5�5�5�5�5�536G6Y6c6�6�6�6�6�6�6�6�6�6�6
7737G7`7q7�7�7�7�7	88+8<8s8�8�8�8�8�8�8�8�899909<9J9[9s9�9�9�9�9�9':8:I:Z:k:|:�:�:�:�: ;	;;&;4;E;Q;_;p;|;�;�;�;�;�;�;<<g<x<�<�<�<�<�<==#=@=I=Z=f=t=�=�=�=�=�=�=�=�=> >1>F>Z>�>�>�>�>�>�>3?G?Y?c?�?�?�?�?�?�?�?�?�?�?   0 �  
0030G0`0q0�0�0�0�0	11+1<1s1�1�1�1�1�1�1�1�122202<2J2[2s2�2�2�2�2�2'383I3Z3k3|3�3�3�3�3 4	44&444E4Q4_4p4|4�4�4�4�4�4�455g5x5�5�5�5�5�566#6@6I6Z6f6t6�6�6�6�6�6�6�6�67 717F7Z7�7�7�7�7�7�738G8Y8c8�8�8�8�8�8�8�8�8�8�8
9939G9`9q9�9�9�9�9	::+:<:s:�:�:�:�:�:�:�:�:;;;0;<;J;[;s;�;�;�;�;�;'<8<I<Z<k<|<�<�<�<�< =	==&=4=E=Q=_=p=|=�=�=�=�=�=�=>>g>x>�>�>�>�>�>??#?@?I?Z?f?t?�?�?�?�?�?�?�?�?   @ �  0 010F0Z0�0�0�0�0�0�031G1Y1c1�1�1�1�1�1�1�1�1�1�1
2232G2`2q2�2�2�2�2	33+3<3s3�3�3�3�3�3�3�3�344404<4J4[4s4�4�4�4�4�4'585I5Z5k5|5�5�5�5�5 6	66&646E6Q6_6p6|6�6�6�6�6�6�677g7x7�7�7�7�7�788#8@8I8Z8f8t8�8�8�8�8�8�8�8�89 919F9Z9�9�9�9�9�9�93:G:Y:c:�:�:�:�:�:�:�:�:�:�:
;;3;G;`;q;�;�;�;�;	<<+<<<s<�<�<�<�<�<�<�<�<===0=<=J=[=s=�=�=�=�=�='>8>I>Z>k>|>�>�>�>�> ?	??&?4?E?Q?_?p?|?�?�?�?�?�?�?   P �  00g0x0�0�0�0�0�011#1@1I1Z1f1t1�1�1�1�1�1�1�1�12 212F2Z2�2�2�2�2�2�233G3Y3c3�3�3�3�3�3�3�3�3�3�3
4434G4`4q4�4�4�4�4	55+5<5s5�5�5�5�5�5�5�5�566606<6J6[6s6�6�6�6�6�6'787I7Z7k7|7�7�7�7�7 8	88&848E8Q8_8p8|8�8�8�8�8�8�899g9x9�9�9�9�9�9::#:@:I:Z:f:t:�:�:�:�:�:�:�:�:; ;1;F;Z;�;�;�;�;�;�;3<G<Y<c<�<�<�<�<�<�<�<�<�<�<
==3=G=`=q=�=�=�=�=	>>+><>s>�>�>�>�>�>�>�>�>???0?<?J?[?s?�?�?�?�?�? ` �  '080I0Z0k0|0�0�0�0�0 1	11&141E1Q1_1p1|1�1�1�1�1�1�122g2x2�2�2�2�2�233#3@3I3Z3f3t3�3�3�3�3�3�3�3�34 414F4Z4�4�4�4�4�4�435G5Y5c5�5�5�5�5�5�5�5�5�5�5
6636G6`6q6�6�6�6�6	77+7<7s7�7�7�7�7�7�7�7�788808<8J8[8s8�8�8�8�8�8'989I9Z9k9|9�9�9�9�9 :	::&:4:E:Q:_:p:|:�:�:�:�:�:�:;;g;x;�;�;�;�;�;<<#<@<I<Z<f<t<�<�<�<�<�<�<�<�<= =1=F=Z=�=�=�=�=�=�=3>G>Y>c>�>�>�>�>�>�>�>�>�>�>
??3?G?`?q?�?�?�?�? p H  	00+0<0s0�0�0�0�0�0�0�0�011101<1J1[1s1�1�1�1�1�1'282I2Z2k2|2�2�2�2�2�2�233$3h3y3�3�3�3�3�3�344$4h4y4�4�4�4�4�4�455$5h5y5�5�5�5�5�5�566$6h6y6�6�6�6�6�6�677$7h7y7�7�7�7�7�7�788$8h8y8�8�8�8�8�8�899$9h9y9�9�9�9�9�9�9
::':k:|:�:�:�:�:�:�:
;;';k;|;�;�;�;�;�;�;
<<'<k<|<�<�<�<`=�=�=�=�=>W>h>s>�>�>%?4?V?   � $  71W1w1�1�1�1�1h2�2323b3s33�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3E4
5*5M5�5�5�7:8i8z8�8�8�8�8�8�89'949S9c9�9�9�9�9�9�9:.:S:c:�:�:�:�:�:;';4;S;c;�;�;�;�;�;�;<<A<Q<v<�<�<�<�<�<=%=J=Z==�=�=�=�=�=>+>M>]>{>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?g?�?�?�?�?�? � D  0#050I0p0�0�0�0�0�0�0�0,1F1\1p1y1�1�1�1�12!2Z2�2�2�2�2�2�2�233=3J3i3v3�3�3�3�3�3�34#4A4R4k4�4�4�4�4�4�4�4�4�4�455!5B5I5V5u5�5�5�5�5�5�5 66)6A6R6k6�6�6�6�6�6�6�6�6�677'7:7N7`7q7�7�7�7�7�7�7�748w8�8�8@:`:�:;.;Q;�;�;�;<<(<4<B<V<<�<�<�<�<�<�<�<�<!=5=G=k=~=�=�=�=�=�=>->A>S>d>y>�>�>�>�>??#?]?}?�?�?�?�?�? � �   0$000>0d00�0�0�0�0�0�0:1K1f1n1�1�1�1�1�122#212`2�2�2333Q3f3�3�4�4�4�4�475X5�5�5�5�5�5�5�5�5	66=6Y6l6�6�6�6�6�6�67707K7\7m7�7�8�8&9F9o9�9�9p:�:�:�;�;<!<H<�<�<Y=|=�=�=�=�=�=?>R>s>�>�>�>�?�? �   0�0T1o1{2�2�2�2�23 3M3a3s3�3�3�3�3�3�34#454F4W4l4�4�4�4�4�4�4�45 515B5w5�5�5�5�5�5�5616C6g6}6�6�6�6�6�6�677$797M7f7w7�7�7�7�7�7�7�78G8V8w8�8�8�8�8 99*9H9b9o9�9�9�9	:-:r:�:�:�:�:�:(;9;�;�;�;G<V<x<�<�<=1=�=�=�=�=�=>*>g>�>�>�>�>�>??:?X?t?�?�? �   70F0P0p0�0�0�0�01'111Q1�1�12&2K2p2{2�2�2�2�2�2�273F3P3p3�3�3�3�3�34?4�4�4�4�45$5F5k5�5�5�5�5�5'666@6`6�6�6�6�6757@7_7�7�7�7�7�7�78'828Q8\8{8�8�8�8�89<9w9�9�9�9�9�9:g:v:�:�:�:�:;!;F;g;�;�;�;�;�;<z<�<�<�<�<=-=8=W=b=�=�=�=�= >\>�>�>�>�>�>?5?�?�?�?�?�?�?   � p   Q0~0�0�0�01W1f1p1�1�1�1�1�12d2�2�2�2(373O3�3�3�3
4/4L4q4�4�4�4�4�4�455h5�5�7�78g8�8�8�8 9;9=U=4?x? � �   ,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�01?1n1�1�1�1B2�2�4�4�56h6P7T7X7\7`7d7h7l7�7�7,8\8�8�8�8�9 :::�:�:�;�;�;�;<<<<< <�<J>�>/?K?�?   � l   (01�1�1�1�2�2�2�2�2�2 3c3�3�4�495i5�5�5�5 7777b7l7�7i8�8�8�8�9�:�:�:�;[<�<�<�<==9=h=�=i>�>N?     |    0$0(0,0004080<0M0�122>3�3g4}4�455a5�5�5�5�5-6�6�7�7�7�7#9.9A9�9�9�95:A:T:�:�:�:;;*;�;�;�;*=?=�=L>|>�>�>�>�?�?    �    00[0u0�0�0$1D1a1�1�1�1�1<2R2f2�2�34444W4�4�45f5�5�5j6r6�6�6:7H7�7�7�7�7#8�9S:�:�:�:�:�;�;G<�=�=�>?4?8?<?@?�?�?     �   00m0�0�0H2I3�3�3�3�3�3 44444444 4$4(4�4�4�45>5^5h5�5�5 6666�6�6�607`7�7�7�78�:�:�:�:�:�:�:�:�:�:;K;|;�;�;�;�;<G<�<=A=M=7>�>�> ??E?�?�? 0 L   0�0!1A1�1�1�12O2n2�2�23o3�3�3`4I5s8�8�8�89W9�9�:%;{;�<�<�=�?�?   @ �   0{0�0�1+2<2t2�2�2�2�2�2�2�2�2�2�2�2�2 3333333t3~3�3.4H4�4�456A78�8>9W:�:�:�:;u;�;@<D<H<L<�<�<�=�>�>�>�>�>?2?�?�?�?�?�?�? P   0#0,0=0[0�0�0�0�0�0�01)1=1O1`1�1�1�1�1�1�12/2@2R2d2�23T3t3�3�3�344+4t4�4�4�4�45)5Q5d5|5�5�56&6�6�6�6�6�6�67"747d7x7�7�7�7�7�78 8D8X8l8�8�8�8�8�89'9t9�9�9�9 ::T:c:�:�:�:
;D;V;�;�;�;�;4<C<q<�<�<�<�<=d=�=�=�=>>#>5>F>R>`>q>�>�>�>�>�>�>�>?J?]?�?�?�?�?�? `    0,0D0�0�0�0
1181[1q1�1�1�1�12%2;2Q2g2}2�2�2�2�2�2�233e3�3�3*4c4t4�4�4�4�4�4�4�4	55#5S5�5�5�5�5�56)6l6�6�6�6�6$737L7f7�7�7�78&8~8�8�8�8�8�8949P9l9�9�9�9�9:':6:N:l:�:�:�:;5;D;Y;y;�;�;�;�;@<G<N<X<l<v<�<�<�<�<�<�<�<�<�<�=�=�=�=a>�>�>p?�?�?�? p 8  40n0u091M1f1�1�1�1�1�12$282Q2e2~2�2�2�2�2 33333333 3$3(3,3034383<3@3D3�3�3#4D4g44�4�4�4�45!545W5o5�5�5�5�5�566A6Y6l6�6�6�6�6�6717I7\77�7�7�7�7�7!8?8R8u8�8�8�8�8�8�89&969K9c9x9�9�9�9�9:+:@:V:f:{:�:�:�:�:�:�:;&;6;K;c;x;�;�;�;�;�;�;<<3<H<^<n<�<�<�<�<2==�=�=�=�=�=>g>v>�>�>�>?&?�?�?�?   � ,  040T0�0�011T1c1�1�1�1
2G2X2{2�2�2�2�2&3k3x3�3�3�3�3<4I4c4�4�455�5�56 696a6{6�6�6�6�6�67787T7n7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7n8�8�8�89929U9m9�9�9�9�9�9:":E:]:p:�:�:�:�:�:;/;M;`;�;�;�;�;�;�;<=<P<s<�<�<�<�<�<=3=K=^=n=�=�=�=�=�=�=>>9>N>f>y>�>�>�>�>??3?H?^?n?�?�?�?�?�?�? � �   00.0>0S0k0�0�0�0�0�0�0�01#1;1�175M5Y5}5-949N9n9�9�9�9:(:E:u:�:�:�:;;\;`;d;h;<<#<E<i<�<�<�<=*=L=s=�=�=�=�=�=�=�=E>�>�>�>?&?E?�?�?   �   (0E0�0�0�01!1N1t1�1�1�1J2l2�2�23f3�34,4�4�4�4�4545R5�5�5�56616A6T6�6�6�6�6�6747Q7d7�7�7�7�7818B8d8u8�8�8�8�8�8�89!929T9t9�9�9�9�9�9:4:L:`:n:}:�:�:�:�:�:�:;C;V;j;y;�;�;�;�;�;<$<D<d<�<�<�<�<==$=6=T=�=�=�=�=�=>4>T>t>�>�>�>�>�>?$?D?d?�?�?�?�?   �   0$0Q0n0�0�011+1N1f1�1�1�12D2]2t2�2�2�2�23"3t3�3�3�3�3�3D4d4�4�4�4�45$5T5t5�5�5�5�56%6<6A6_6�6�6�67$7d7�7�7�7
8,8N8l8�8�8909T9t9�9�9:4:T:q:�:�:�:�:�:;;!;4;T;k;;�;�;�;�;�;!<1<D<[<o<}<�<�<�<�<�<=!=4=d=�=�=�=�=>$>D>d>�>�>�>�>?4?d?�?�?�?�?   �    0$0D0d0�0�0�0�0111T1t1�1�1�1�1242T2t2�2�2�2�2343T3t3�3�3�3�3444T4t4�4�4�45545T5t5�5�5�5�5�5�566D6Q6d6�6�6�6�67$7D7d7�7�7�7�788D8d8�8�8�8�899/9=9L9^9�9�9�9�9�9�9(:M:c:z:�:�:�:�:�:�:;1;E;S;b;t;�;�;�;�;<(<8<d<�<�<�<�<==D=d=�=�=�=�=�=>4>Q>t>�>�>?$?D?d?�?�?�?�?�?   � �   040T0q0�0�0�0$1I1l1�1�1�12242Q2d2�2�2�2�2�23!343Q3a3t3�3�3�3�3444^4�4�4�4�4�4515N5t5�5�5�5�56(6;6�7�7�7�7�7�7�7�7�7�7�7�7�7�7888�8�8�8X9k:}:�:�:�:�:�:�:;D;d;�;�;�;<D<d<�<�<�<�<�<=4=Q=a=q=�=�=�=�=>1>W>�>�>�>�>�>?4?g?�?�?�? � �   0T0g0{0�0�01!1A1a1�1�1�1�12H2Y2�2�2�2�233F3P3�344k4�4�4�45!545h6�6�6�6Y7^7�7'9T9q9�9�9�9�;�;�;<�<�<^>�>�>�>�>�>??1?[?�?�?�? � �   030;0A0F0s0�0�0191a1�1�1�1�1�12<2C2r2�2�23/3�3-4a4{4�4�4o5�5�56D6q6�6�6�6�6777d7�7�7�7�78"868[8o8�8�8�8�8949S9s9�9�9�9�9�9::>:R:f:�:�:�:�:�:;7;g;�;�;<T<t<�<�<�<=7=a=�=�=�=>4>T>�>�>�>?*?W?�?�?�?   �   070i0�0�0�0<1w1�1�1�1�1�12�2�23�34K4m4�4�4�4515Q5�5�5�56D6a6�6�6H7`7z7�7�7�7�78/8A8�8�8�8�89'9`9}9�9�9�9|:�:�:�:;�;�; <@<�<�<�<=,=B=n=�=�=�=�=">4>�>�>?k?�?�?  �   0B0�0�0�0+1a1�1�1�12?2{2�2�273�3G4s4{4�4�45>5�5�56,6N6b6t6�6�6�6+7j7�7�7	8V8x8�8�89!9Y9t9�9�9:::t:�:�:�:;<;P;�;�;�;q=y=�=�=>�>?,?I?r?�?�?     �   0Q0�0�0�0141t1�1�1�1D2�2�2D3�3�344�4�4$5t5�56d6�67Q7�7�748t8�89k9�9�9T:�:�:;K;�;�;�;$<[<�<�<�<=^=�=�=A>a>z>�>�>�>'?W?�?�? 0 �   0O0�0�01D1n1�1�1�1$2T2�2�2�213d3�3�3414g4�4�4�4Q5�5�5�5�56Q6e6x6�6�6�67!7t7�7�7�7�7�7 8888A8u8�89$9Y9�9U:�:(;,;0;4;8;<;@;D;H;p;B<�<�<�<�<�<�<�<�<�<�=�=�=�=�=�=�=8>�>�>�>�>�>�>$?P?   @ �   070!1d1�1F2t2�2�2�23$383H3w3�3�3�3�3�3 44,4@4]4k4}4�4�4�4�4�4$5D5d5�5�56616P6a6�6�6�6�67/7B7�7�7�7�7B8W8h8t8�8�8�8�89989L9^9o9�9�9�9�9�9�9:,:l:�:�:�:�:;J;k;�;�;�;V<�<�<�<=$=)=>=m=�=�=�=�=R>d>�>�>?9?�?�?�?�?�?�?   P �   00,0=0P0l0�0�0�0!141V1�1�12g2�2353�3I4k455�5�5�5�6�67#7�8�8�89$9T9t9�9�9�9�9:4:Q:n:�:;5;S;�;�;�;�;=<I<h<�<�<�<N=Z=y=�=�=
>)>]>�>�>�>?�?   ` �   e01l1}1�1�1�122c2k2{2�2�23#3G3O3�3�3�34#4+4�4�4�4�4�4
5.5k5�5�5�5�5&6Q6�6�6�6�6�6777Q7[7c7p7~7�7�7�7�7�7�7�78}8�8�8�8�8�8�8 999P9w9�9�9�9�9�9�9�9�9:::#:1:I:�:�:;�;�<*=z=W>�?�? p �   "0�0 111111�1�2<3F3�3�3�3R4�4�45)5�56U6�67Z7�7�7�7�7!8F8Z8�8�8+9?9�9�9::|:�:�:$;(;,;0;4;8;�<==V=^=f=n=�=�=�=�=�=\>�>�>�>�>�>�>�>"?N?�?�?�?   � �   i0y0�0�0�0�0'1Q1b1�1�1D2H2L2P2T2a2t2�2�2�23G3�3�3�3'4W4�4�4�45!5D5w5
6=6W6�6�6�6$7D7d7�7�7�7�8�8�8�8�8949M9z9�9�9�9:1:D:t:�:�:�:;1;T;�;�;�;<!<A<a<�<�<�<�<=4=T=t=�=�=�=�=>$>D>d>�>�>�>�>�?�? � |   0�0�0F1g1�1�1'2�2323�3@4Z4�4M5i5�5�5�5<6�6�6�6	7G7�7�78�8�8�8�879�9:9:T:i:�:;�;�;!<�<�<�<�<'=�=>*>�> ?:?�?�?   � �   040T0t0�0�0�0"1S1r1�1�1�1�12/2=2�2�2�2�23$3A3T3�3�3�3�3'4T4�4�4�4�4�4545T5t5�5�5�5�5�5�566$6D6d6�6�6�6�67D7d7�7�7�7/8g8�8�8949Q9a9�9�9:$:W:�:�:�:�:$;A;d;�;�;�;<4<T<�<�<�<�<=$=D=W=q=�=�=�=�=�=>$>G>t>�>�>�>�>�>�>�>?%?6?T?t?�?�?�?�?�? � �   0"020T0t0�0�0�0�0141Q1d1�1�1�1�1�12$2D2d2�2�2�2�2313P3q3�3�3�34D4d4�4�4�4�45!545T5t5�5�5�5�56646Q6e6u6�6�6�67W7�7�7�7�7848T8t8�8�8�89$9J9|9�9�9�9�96:g:�:�:�:!;G;q;�;�;�;�;6<S<z<�<�<�<=$=D=d=�=�=�=�=>>D>l>�>�>�>�>�>$?<?e?}?�?�?�?�? � �    00D0\0�0�0�0�0�01 101d1�1�1�1�1�12D2m2�2�2�2�2�2$3D3d3�3�3�3�3444T4q4�4�4�4�4�45!545t5�5�5�5�5646T6t6�6�6�6�67747T7t7�7�7�78$8Q8t8�8�8�8949Q9t9�9�9�9�9:D:q:�:�:;D;t;�;�;�;0<O<g<�<�<�<=!=D=T=�=�=�=�=>2>U>s>�>�>�>
??7?[?l?�?�?�?   � �   010Q0q0�0�0�0141T1�1�1�1272a2�2�2�2�2343d3�3�3�3	4'4D4q4�4�4�4�45D5w5�5�5�556O6�677o7�7�7�7�78;8j8�8�89$9T9�9�9�9�9:$:A:d:�:�:�:;$;A;d;�;�;�;�;$<Q<t<�<�<�<�<=1=@=d=�=>$>W>�>�>�>?a?�?�?�?   � �   040i0�0�0�0�0�01�1�172D2�2�2�2 3�417J7�7�7�7�7%8g8�8�9�9�9�9:4:T:|:�:�:�:B;U;Z;t;�;�;�;D<d<�<�<�<�=�=�=>'>g>�>�>�>?;?@?�?�?�?�? � �   010T0t0�0�0�01$1A1d1�1�1�1O2�2�2�2�3444%4,434:4A4H4�4555�5G6%717X7]7�7818T8q8�8�8�89$9U9a9t9}9�9�9�9�9:D:q:�:�:�:;$;D;�;�;�;`<�<�<#=[=�=�=�=5>:>e>s>>�>�>�>�>�>�>??2?]?w?�?�?�?�?�?�?   4  00+070E0g0x0�0�0�0�0�01$151U1o1�1�1�1�1�1�1�1
22'252W2h2�2�2�2�2�2�23%3E3_3p3|3�3�3�3�3�344E4T4`4r4�4�4�4�4�4�4�45=5W5h5t5�5�5�5�5�5 666<6M6m6�6�6�6�6�6�67707C7j7�7�78.8�8�8�8�8�89,9@9`9t9�9�9�9�9E:V:a:o:�:�:�:;%;9;K;\;�;�;�;�;!<2<;<D<V<a<{<�=�=�=�=�=�=	>>>'>1>?�?�?�?�?�?�?�?�?�?    �   �1�1�1(2U2k2)30373>3E3L3S3Z3a3h3o3v3B4u4�4�4�4U5y5�5�5656]6�6�6�67U7�7�7�78E8�8�89B9g9�9�9�91:Y:�:�:�:�:�:;1;Y;�;�;�;7<f<�<�<=M=�=�=>B>u>�>�>2?e?�?�?   �   50u0�0�0%1U1�1�12b2�2�2363p3�34E4�4�45U5�5�5$6X6s6�6�6�6�67B7�7�7�7(8�8�8%9h9�9�9�9%:h:�:�:;U;�;�;<R<�<�<=D=�=�=>T>Q?�?�?�? 0 �   80�0�0%1e1�1�1%2e2�2�2%3r3�3�3424e4�45E5�5�56�67u7�7�768b8p8t8z8~8�8�8�8�859u9�9�95:�:�:d;�;�;�;<7<R<~<�<�<=,=E=s=�=�=>1>d>�>�>�>?J?�?�? @ �   *0?0~0�0�0�0J1m1�1�1�1�1�182j2�2�2�2�2$3t3424h4�4�4�4�4555u5�5�56U6�6�6%7e7�78B8�8�89U9�9�9:$:1:7:f:m:�:�:�:�:;;;;;;,;4;W;<<"<e<t<�<I>�>�>�?   P �   0�2�273<3|3�3d4�4545d5�5�5�5�5;6G6�6�677.797Q7�7�7�7�7�788*8D8l88�8�8�8�8�8�8a9�9�9�9�9:1:T:d:�:�:�:�:;4;a;�;�;�;�;<!<D<d<�<�<�<�<!=A=d=�=�=�=4>t>�>�>?4?T?t?�?�?�?   ` <   0$0A0d0�0�0�0:1a1�1O9T9�9�9X:]:�:�:^;j;�;�;�;�;�>�> p 4   �4h5l5p5t5x5�798D8L8^84;�=�=5>u>�>�>5?u?�?�? � �   0U0�0�01E1�1�1�1"2R2�2�2�253u3�3�354u4�45U5�5�556u6�6d7�7�7M8a8k8�8�8z9�9�9�9�9%:-:P:h:;';;;K;W;`;�;�;�;�;h<p<x<�<�<�<�<>>#>+>�>�>�>�>�>�>�>
?/?M?Y?e?q?}?�?�?�?�?�?�? � �   0000A0J0b0n0z0�0�0�0�0�011�1�1�1�1222A2�2�23n3v3~3�3�3�3�34#4�4g5z5�5�5�5@6H6y6�6�6�6�6�6�677.7:7P7Y7b7�78K8_8�8�8�8�89!9�9,:=:m:u:�:�:�:#;,;7;z;�;<J<V<�<�<=U=a=�=>@>�>�>??/?r?   � �   �0�0�0�0�1�1�1�1222A2�2�2�233B4�4�4'5<5E5N5b5�5�5G6a6j6r6�6�6�6�8�8�8�8�8�8�8�8979U9\9`9d9h9l9p9t9x9�9�9�9�9�9::E:`:g:l:p:t:�:�:�:�:�: ;;;;;;^;d;h;l;p;�<=s=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>O>T>^>�>�>�>�>�>?;?V?�?�?�? � �   >0l0�0�01#1B1Y1h1�1�1
222|2�2�2�2�2@3Q3�3�3�3�3�3�3G4S4[4�4�4�45C5K5S5�5�6�6�6q7y7�7�7�7�78818=8I8�8�8�8�8�89�9�9�9�9+:2:::�:�:�:�:�:�:	;";Y;i;K<�<�<�<�=�=o>v>�>�>�>�?�?�?�? � �   '0<0c0�3�466>6D6c6i68.:2:6:::>:B:F:J:D;x;�;�;�;�;�;<<%<+<1<7<><E<L<S<Z<a<h<p<x<�<�<�<�<�<�<�<�<�<�<�<=Q=�=Z>j>v>�>�>�>�?   � �   0�0,1O1]1t11�122$2>2]2r2|2�2�2�2�2�2�2�2�2U3�3�3�3�3�3�3494E4Q4g4�4�4�4�4�4�4�4�4�4�45'505s5w5{55�5�5�5�5�5�5�5�5�5�5�5�5u6�6�6�6�67B7�7�7�7�7�78"8b8�8�8�8�8!9,9>9R9�9�9�9�9":�:�:�:;�;4<R<r<�<='=9=D=q=|=�=�=�=2>=>O>b>x>�>O?�? � 4   o1�1�1�67V79�9�<�<�<=>�>�>"?*?s?�?�?�?�?   � �  0#0/0>0c0�0�0 1"1=1V1g1{1�1�1�1�1�1�1�1�1�1�12'2-282F2O2Y2i2n2s2�2�2�2�2�2�2�2�2333$343@3E3P3Z3p3�314H4U4a4q4w4�4�4�4�4�4�4�4 55505_5f5t5}5�5�5�566O6n6�6�67	77e7�7�7818Q8w8�8�8�8�8�8�89!9�:�:�:;G;S;_;n;y;�;�;�;�;�;�;<"<3<g<�<�<�<�<�<�<�<�<�<�< ====1=;=A=\=l=u=}=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>
>>>>%>*>0>8>=>C>K>P>V>^>c>i>q>v>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?	????!?'?/?4?:?B?G?M?U?Z?`?h?m?s?{?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?        00
0000&0,0:0H0O0\0e0�0�0�0�0101G1L1g1l1�1�12�2�2�2�23�3�3�3�3�344]4u44�4�4�4�4�4�4�4�4�4�45!5O5b5�5P6�6�6S7e7�7�7�7�7�7"8�8�8�8�899 9:":*:0:<:A:F:K:T:�:�:�:�:�:�:;;;v;�;�;�;<�<�<�<�<�<"=�=�=�=�=�=�=�= >>>&>1>9>F>P>v>�>�>�>�>?V?j?�?�?�?    �   0�0�0}1�1�1�1T2!3P3Y3�3�3�4�4�4�4�5�5�6�6�7�7�78h8�8�89<9[9::::T:�:@;�;-<�<'===v=�=�=>,>3>:>A>Y>h>r>>�>�>�>?9?     �   �0�0�011$1O1�1�12!2,2C2]2x2�2�2�2�2�2�223h3{34?4f4�4�5�5�6�6�7�8�8�8�8D9Q9}9�9�9�9t:�:�:�:�:�:I;U;];i;�;�;�;<<6<X<�=�=�=�=�>�?�?�?�?�?�?   0 �   *020F0P0n0z0�0�0�0�0�0�0 111$101d1n1v1�1�1�1�1�1�1222T2c2k2q2�2�2�2�2�2)353E3Q3n3t3�3�3�3�3~4�4�4�4�45*5K5o5{5�5�6�677H7�7�7A8x8�8�8�89�9�9�9�9�9:!:7:@:K:S:q:}:�:�:�:�:T;�;�;�;�;<<D<d<�<~=�=�=�=&>.>T>x>�>�>�>�>[?�?�? @ h   0&0H0�0	181w12#2;2C2d2�2�3
444�4X5�5�5&6E6�6�6�6�6�6�6�67c7o7�7 88�8�8�9�9�9::;�=�>�>   P �   �0�0�0�0T1f1x12)2/292O2b2x2�2�2�2�2�2363;3`3u3{3�3�3�495D5�6�67)7�8�8999 9$9(9Q9w9�9�9�9�9�9�9�9�9�9:::::z:�:�:�:�:�:�:�:�:1;8;<;@;D;H;L;P;T;�;�;�;�;�;&=?�? ` �    1v3{3�3�3�3�3d4�4�4�4�4\5b5n5�5�5	666�78
8.8=8`8q8w8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999.9F9L9U9[9e9p9�9�9�92:::F:�:�:�:�:;u;�;�;�;�;<<<�<�<�<=='=c=�=�=�=�=???�?�?�?�?   p �   00y0�0�0�0�0121:1W1g1s1�1?2`2g2�2�2�2�2�3�3�3�354s4�4�4�45"555W5^5�5�566�6�6#727Q7�7�7�7�7�7	88-8?8Q8c8u8�8�8�8�8�8�8�<�<i=X>�>
?�?�? � X   �011�1�1�1�2�2�2�2�2�2X3z4�4*6�6�6V7^7j7y788S8�8�9�9�;.<:<�<�<�<�<w=�=�=P>   � 4   �1�165:5>5B5F5J5N5R5V5Z5^5b5p5.6G6V6w6�67   � D   H1�3b4�4�4�4�4�4I5Z5n5t5y5a7�7�7�7N8�8�8�8R9X9b9k9t9�9�9�9   � �  �011111$1(1,1P2T2X2\2`2d2h2l2p2t23 3$3(3,3034383<3@3D3H3L3P3T3X3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;===== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � d   00000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; � @  @3D3H3L3P3T3X3\3`3d3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444 4$4(4,4044484H4L4P4T4X4\4`4d4h4l4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555555054585<5@5D5H5L5P5T5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666 6$6(6,60646D6H6L6P6T6X6\6`6d6h6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 888 8$8(8,8084888<8P8T8X8\8`8d8h8l8p8t8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 94989<9@9D9H9L9P9T9X9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::: :$:(:,:0:4:8:<:P:T:X:\:`:d:h:l:p:t:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;;; ;$;(;,;@;D;H;L;P;T;X;\;`;d;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<(<,<0<4<8<<<@<D<H<L<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<=== =$=(=,=0=4=8=L=P=T=X=\=`=d=h=l=p=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$><>@>D>H>L>P>T>X>\>`>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ?????(?,?0?4?8?<?@?D?H?L?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � �  0000 0$0(0,00040�0�0�0�0�0�0�0�0�0�0(1,1014181<1@1D1H1L1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 222 2$2(2,2024282<2T2X2\2`2d2h2l2p2t2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2333333 3$3(3,3\3`3d3h3l3p3t3x3|3�3�3�3�5�5�5�5�5�5�5�5�5�5�5(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8   � <  p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�1�1 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,303L4P4T4X4\4�4�4�4�4�4�4555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5�5�5�5�5�5�566�6�6�6�6�6�6�6�6 77777777 `    �0�0�0   �    $2(2 � 8   ?$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?   � �  �9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;$;,;4;<;D;L;T;\;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? �   0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88 �    �:�:�:�: �    
6666 0 �   p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9   ` $  ::�:�:�:�:�:�:�:�:�:�:�:�:;;,;0;@;D;H;P;h;x;|;�;�;�;�;�;�;�;�;�;�;�;�;<<<< <8<H<L<P<X<p<�<�<�<�<�<�<�<�<�<�<�< ====,=0=4=8=<=D=\=l=p=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>,>0>4>8>L>P>`>d>h>l>p>x>�>�>�>�>�>�>�>�>�>�>�>??????4?D?H?X?\?`?d?h?p?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   p d   00(0,0<0@0D0H0L0T0l0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01$1(181<1@1D1H1P1h1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12 2$24282<2@2D2L2d2t2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233 3034383<3@3H3`3p3t3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3444,4044484<4D4\4l4p4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4555(5,5054585@5X5h5l5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 666$6(6,60646<6T6d6h6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�677 7$7(7,70787P7`7d7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7888 8$8(8,848L8\8`8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�89999 9$9(909H9X9\9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9 ::::: :$:,:D:T:X:h:l:p:t:x:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;; ;(;@;P;T;d;h;l;p;t;|;�;�;�;�;�;�;�;�;�;�;�;<<<<<4<D<H<X<\<`<d<l<�<�<�<�<�<�<�<�<�<�<�<�<�< ===$=4=8=H=L=P=T=\=t=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>$>(>8><>@>D>L>d>t>x>�>�>�>�>�>�>�>�>�>�>�>�>�>???(?,?0?4?<?T?d?h?x?|?�?�?�?�?�?�?�?�?�?�?�?�?   � H  0000 0$0,0D0T0X0h0l0p0t0|0�0�0�0�0�0�0�0�0�0�0�01111141D1H1X1\1`1d1l1�1�1�1�1�1�1�1�1�1�1�1�1�1 222$24282H2L2P2T2\2t2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23$3(383<3@3D3L3d3t3x3�3�3�3�3�3�3�3�3�3�3�3�3�3444(4,40444<4T4d4h4x4|4�4�4�4�4�4�4�4�4�4�4�4�45555 5$5,5D5T5X5h5l5p5t5|5�5�5�5�5�5�5�5�5�5�5�56666646D6H6X6\6`6d6l6�6�6�6�6�6�6�6�6�6�6�6�6�6 777$74787H7L7P7T7\7t7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78$8(888<8@8D8L8d8t8x8�8�8�8�8�8�8�8�8�8�8�8�8�8999(9,90949<9T9d9h9x9|9�9�9�9�9�9�9�9�9�9�9�9�9:::: :$:,:D:T:X:h:l:p:t:|:�:�:�:�:�:�:�:�:�:�:�:;;;;;4;D;H;X;\;`;d;l;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<$<4<8<H<L<P<T<\<t<�<�<�<�<�<�<�<�<�<�<�<�<�< ===$=(=,=0=4=<=T=d=h=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>> >$>(>,>0>8>P>`>d>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>??? ?$?(?,?4?L?\?`?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?   � t  0000 0$0(000H0X0\0l0p0t0|0�0�0�0�0�0�0�0�0�0�01111101@1D1T1X1\1d1|1�1�1�1�1�1�1�1�1�1�1�1�1�1 22242D2H2\2`2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2 3333(3,3<3@3D3L3d3t3x3�3�3�3�3�3�3�3�3�3�34444 4(4@4P4T4d4h4p4�4�4�4�4�4�4�4�4�4�4�4�455505@5D5T5X5`5x5�5�5�5�5�5�5�5�5�5�5�5�566 60646<6T6�6�6�6�6�67$7@7L7h7�7�7�7�78(8H8d8h8�8�8�8�8�8�89909P9p9�9�9 � P  $0(02222 2$2(2,20242�2�2T9X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<$<D<P<T<X<\<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=�>�>�>�>�>�>�>�>�>�>�>?????? ?$?,?0?P? � �   X2p2�2�2�2�2�23,3D3`3|3�3�3�3�34(4D4`4|4�4�4�4�45(5D5`5|5�5�5�5�5606L6h6�6�6�6�6�6787X7t7�7�7�7�78 8@8`8�8�8�8�8 9 9D9h9�9�9�9�9:<:\:|:�:�:�:;@;h;�;�;�;<@<h<�<�<�<=<=l=�=�=�=>H>t>�>�>�> ?L?x?�?�?   � T   0,0X0�0�0�0101X1�1�1�1242`2�2�2�23<3`3�3�3�3�34,4H4d4|4�4�4�4�4505P5t5                                                                                                                                                                                                            