MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��Ƿڵ��ڵ��ڵ�)zr��ڵ���T��ڵ���j��ڵ���U��ڵ�j%~��ڵ��ڴ��ڵ���T��ڵ���i��ڵ���k��ڵ�Rich�ڵ�                PE  L ��DT        � !  �  �     �     �                         �	         @                   �� K   ̚ (                             	 �{  @� 8                           0l @            � �                           .text   %�     �                   `.rdata  `�  �  �  �             @  @.data   E   �  &   �             @  �.reloc  �{    	  |   �             @  B                                                                                                                                                                                                                                                                                                                                                                                        hС衩 Y�������������������������������������U��D���D� P���V=�  v3�^��]�jhh�h�   j���    �2� ����t���ı ����
���    jhh�h�   j� � ����t��蒱 ����
���    輵 ����M�D����    Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M���(�@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�ЍE�P�u� �D��M�Q�@�@�Ѓ����D�V�@�@�СD��M�VQ�@�@�Ѓ��C  �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�$�TF  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ���F  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ��n  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ���W  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ��@^  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ��{_  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ��&a  ��ul�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�Ѓ��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��MЃ��@Q�M��@x�ЋD�����E�P�I�I�у���tZ�D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��M���Q�M�QP��  ���A  �D��M�Q�@�@�Ѓ��>  �M��@� �D��M�jh�  �@�@4�СD��M�jh�  �@�@4�СD��M�jWh�  �@�@4��j�E�Ph&� �+� ���M��@� �D��M�Q�@�@�СD��M�Q�@�@�Ѓ��   ^��]��V�5����t����� V蘄 ���5�����    ��t���ګ V�t� �����    ^������U��D���   �SP���VW=�  v	3�_^[��]ËE=�  ��  t#�� ��  Hu۹���!� �����_^[��]Ë��   ���   ��jjP�E��i� ���M��ު �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@Qj�M��@8�СD��M�Q�@�@�СD����M����   ���   �Ѕ���  �E��� ��	 �
��$    �I �D��M����   ��?���P���   �ЋD��؋��   �ˋRx�ҋD����E�P�I�I�ыD��A�M�QV�@�Ѓ����� �ˉE�賀 �    t�D��M�Q�@�@�Ѓ���  �Eԋ�P��p���P葀 ��躇 ��p���蟅 �D��Mԋ@�@<�Ѕ�uT�D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�M�Q�@�@�СD��M�Q�@�@�Ѓ� �D�����@V�@�СD��M�VQ�@�@�Ѓ��E�P�#  �ȃ���tL�D��U�RW�@�@8�СD��M�Q���W�@�@8�СD��u�����P��'  P�B4���   �M�詨 �D��M�Qj�M��@�@8�СD��M�QW�M��@�@8�СD��M�Q���W�@�@8�СD��u�����P��'  P�B4�СD��M��]�QS�@�M��@D��C�M��]�腨 �D��M�Q�@�@�СD��M�Q�@�@�Ѓ��D�G�M����   ���   �Ѝ�?���;�������D��M�Q���h�	 �@�@D�ЍM��� �D��M�Q���   ���   �Ѓ��   _^[��]�=�  �F����[  j �jM  ���"M  _^�   [��]�������U���M�\M�YM�XM�M�E]����������������U���EW�f/�v
�M�E]����f/�w��E�E]��������������U���UW�f/����v(��	f/�v(��]f/�v(��	f/�v(��ef/�wf/�v�E(�� �X�P]�(ċE� �X�P]����U���E�Mf/�v
�M�E]��E�E]����������U���E�Mf/�v
�E�E]��M�E]����������U���E�M4f/�w(��M�U,f/�w(��U�]$f/�w(ӋE��H�@]��U����E���Vd ����]��E��\�fTP��\��M��E���]�U���E��f/���E�$v
� � ��]��� ��]��U���M�\M�YM�XM�M�E]����������������U���M$�\M�U<�E�Y��XM��M,�\M�Y��XM�H�M4�\M�Y��XM�H]�������������U���E�\Ef.���E���Dz��]��E�e�u]��U���E�M�Y���Y���X��E�Y@��X��M�E]�����U���E�XE�XE�Y���E�E]�������������U���M�Ef/�v(��E�Mf/�v�M�E]�U���E�M�Y���Y`��X��E�Y0��X��M�E]�����U��EP�u�` �E��]����������U��EP�u�a �E��]����������U���MW��U�\�f.ȟ��D{�E�\��^��E�E]������������U���MW��e�\�f.ȟ��Dzf(���U,�\��^�f.ȟ��Dzf(���]$�\��^�f.ȟ��D{�E�\��^��E� �X�P]���������U���M�\M�YM�XM�M�E]����������������U���M�UE�Ef��\�f�fY��YU,fX��X� �P]������U���M���f.ʟ��Dz�E]�W�f/�r��]��]f/�s��^�(�(��:n �E�E]�U��������U$f.ӟ��Dz�E�oE� �~Ef�@��]�W�f/�r�M��1�Ef/��E�s!(��^���m �U$W�����E�f/�r�M��)�Ef/��E�s(��^��m �U$W��E�f/�s(f(��Mf/�sf(�����^��Xm f(ȋE�E��@�E���@��]������U����eW�f.��E����Dz�E��]����f(��^�f.ӟ��Dz�E�E��7f/�s1�Mf/��M�s!(�(��^���l ����e�E��E�\�f(��l �YE��E�E��]�������������U����]W����f.��E���Dz�U�U��   f(��^�f.���Dz�E,�E��4f/�s)�U,f/��U�s�^�(��l ����]�E��E�\���k ���f(��Ye�W��]�U�e�f.؟��Dz�U��{f(��^�f.���Dz�E$�E��4f/�s)�U$f/��U�s�^�(��xk ����]�E��E�\��Xk �]f(��YM�W��U�M�f.؟��D{x���f(��^�f.���Dz�E�E��7f/�s1�Mf/��M�s!(�(��^���j ����]�E��E�\�f(���j f(��YU��E�E��@�E���@��]�������������U���E�Mf/�v
�M�E]��E�E]����������U���M4�Ef/�w(��U,�Mf/�w(��]$�Uf/�w(ӋE��H�@]��U���E�M]������U���E�YE$�E� �E�YE,�@�E�YE4�@]�������������U���Uf.�����Dz��]����f(��\E�^��\��M�E]����U���]W����f.ٟ��Dz(��f(��\E4�^�(��\��ef.���Dz(��f(��\E,�^�(��\��mf.���D{f(�(��\E$�^��\ȋE��`�X]�������������U���E�XE���f/�vW��E�E]��\��E�E]�����������U���EW��XE4���f/�v(���\��M�XM,f/�v(���\��e�Xe$f/�w(��\ڋE��H�@]�������U���U�E$�XU�XE,�]�e4�E�X��X��Y���Y��f/�v�oE� f�X]��oE$� f�`]���������������U���E�Mf/�v
�E�E]��M�E]����������U���E�M4f/�w(��M�U,f/�w(��U�]$f/�w(ӋE��H�@]��U�����f(�f(��\M�\E�Y��\��U�E]��U������Ef(��\Mf(��\E$�Y�f(��\�f(��\M� f(��\E,�Y�f(��\�f(��\M�@f(��\E4�Y��\��P]�������������U���E���f.����DzW��E�E]��\��E�^��E�E]���U���]W����f.ٟ��Dz(��f(��\��]4�^��ef.���Dz(��f(��\��e,�^��Ef.����D{�U$�\��^ыE��`�X]����������U���E�E]������U���E�XE$�E� �E�XE,�@�E�XE4�@]�������������U���U�E$�XU�XE,�]�e4�E�X��X��Y���Y��f/�v�oE� f�X]��oE$� f�`]���������������U������]f/�v
�E�M��]����f(�(��\M�\��Y��Y��\��U�E]���������������U���5���e4f/�����-�v�]�Y��Y��!f(�f(��\M�\�f(��Y��Y��\��},f/�v�e�Y��Y�� f(�f(��\M�\�(��Y��Y��\��}$f/�v �U�E�Y��`�X�Y��]ËEf(��\Mf(��\��`�X�Y��Y��\��]������U����������ef/�vC�M(��Y�����\�(��Y��Y��Y��Y��X��$�$��]��E�p �M�Y�����\��\]�Y��M�Y��Y��X��$�$��]�����U�����m4�����f/�v9�%�(�����Mf(��Y��\�(��Y��Y��Y��Y��E�E��o �%�f(��M4����E�Y��Y��\��Y�f(��\M4�Y��m,�X����f/��\$v)�M(��Y�f(��\�(��Y��Y��Y��Y��E�E�Vo �%�f(��M,����E�Y��Y��\��Y�f(��\M,�Y�����X��$�]$f/�v)�M(��Y��\�(��Y��Y��Y��Y��X��A�E��n �M$�Y�����\��\U$�Y��M�Y��Y��XЋE�$�@�D$��@��]������U������Uf/��]v@W�f.؟��Dz
�E�E]��Y����(��\��^��\��M�E]����f.؟��DzW��E�E]��\��\��Y��^��U�E]���������U���-��W��U4f/��=��]�%��v(f.ٟ��Dz(��<�Y�f(��\�(��^��\��#f.ܟ��Dz(���\�f(��\��Y��^��],f/��uv(f.���Dz(��<�Y�f(��\�(��^��\��#f.����Dz(���\�f(��\��Y��^��u$f/�v9�mf.���D{L�Y�f(ċE(��\��X�P�^��\��]��Ef.ğ��D{(��\��\��Y��^̋E��X�P]����U������Ef/�v6�Y�����XEf/�vW��E�E]��\��E�E]��\��Y��XE�E�E]����������U�����W��E4f/��5���-�v�Y��XEf/�v(���\���\��Y��XE�M,f/�v�Y��XMf/�v(���\���\��Y��XM�e$f/�v)�Y��Xef/�w*�E(��\��H�@�]�(��\��Y��XU�E��H�@]��������U������Ef/�v'�Y��Mf/�v
�M�E]��E�E]��\��M�Y�f/�v
�M�E]��E�E]���������U������E4f/����]v
�Y�f/���\��Y�f/�w(��E,f/��ev
�Y�f/���\��Y�f/�w(��E$f/�v�M�Y�f/���\��M�Y�f/�w(ȋE��`�X]�����U���%��W��Mf/��m���v,f.���Dz(��?�Y�f(��\�(��^��\��"f.���D{(�\�f(��\��Y��^�f/�w
�U�E]��]�E]���U���%�����M4W�f/��-��u���v(f.���Dz(��7�Y�f(��\�(��^��\��f.���D{!�\�f(��\��Y��^�f/�w�U���]��M,f/��uv(f.���Dz(��7�Y�f(��\�(��^��\��f.���D{ �\�f(��\��Y��^�f/�wf(��f(��M$f/��uv(f.���Dz(��7�Y�f(��\�(��^��\��f.���D{�\�f(��\��Y��^�f/�v(ӋE�E���x�@��]���������U���E�\EfTP��E�E]��U���E�\E$�E�P�fT�� �E�\E,fT��@�E�\E4fT��@]���������U���Mf(��Y��XU�YM�\��U�E]�����U���M��f(��XU$�E�Y��YM$�\��M�f(��XU,�Y��YM,�\��M�Pf(��XU4�Y��YM4�\��P]��U���E�e]������U���E$�\E�E� �E,�\E�@�E4�\E�@]�������������U���EW�f/��Uvf/�v
�M�E]��^��E�E]�������������U���MW�f/��U4vf/�v(���^��Uf/��],vf/�v(���^��ef/��]$vf/�w(��^ËE� �P�H]�������������U���H�oE�E�P�E�E��~EPf�E��H �oE$�E�P�E�E��~E4Pf�E��H �U��E��E��M�P�uf��U�f�M��J �E����]������U���H�oE�E�P�E�E��~EPf�E��)H �oE$�E�P�E�E��~E4Pf�E��H �UЍE��E��M�P�uf��U�f�M��I �E����]������U���H�oE�E�P�E�E��~EPf�E��G �oE$�E�P�E�E��~E4Pf�E��G �UЍE��E��M�P�uf��U�f�M��I �E����]������U���H�oE�E�P�E�E��~EPf�E��)G �oE$�E�P�E�E��~E4Pf�E��G �UЍE��E��M�P�uf��U�f�M��H �E����]������U���U�E$�XU�XE,�XU�XE4�Y���Y��f/�v�E���f� �@]ËEW�f� �@]�������������U���M$�U,�]4�\M�\U�\]����E�X��X��X���P�X]���������U���M$�U,�]4�XM�XU�X]����E�\��\��\���P�X]���������U��E �� H��   HtuHt;�E�M�Y���Y`��X��E�Y0��X��M��E���]��oE�~U(�f�f/��E�w�M�f/�vbf(��M��E���]��E�XE�XE�Y���E��E���]��E�M�Y���Y���X��E�Y@��X��M��E���]�����������U����u,�oe���]$��� f�X������M���E�E�]��U��\��\��\��Y��Y��Y��X��X��X�f�� f�X��]��������������U���MW�f/�v��]���f/�r�^X��M�E]��X(��^��(�����S �E�E]��U���MW��X���f/��%(��-���5�v�E��T��f/�r�^��M��;�X��^�(�(��iS �X��%(��-���5��E�W��Mf/�v(��6��f/�r�^��"�X��^�(�(��
S �X�f(�W��Uf/��M�w<��f/�r	(��^��%�X(����^��(��R �M��E� �E��H�@��]������U���MW���f/�r�M��E���]�(�����`R �E��E���]�����U����MW�f/�����M�s(�(��$R ����E�W��Uf/��U�s(�f(���Q �E�W��Mf/�s(������Q f(ȋE�E��@�E���@��]���U��D��MQ�@�@�Ѓ�]��������U��D���4�@S�]��V�@`Wj �Ћ�   �����   �I V��訆 =�   ��   �D���V�@�@T�Ћ��MܡD�Q�u��@�@�СD��M܃��@Qj�M̋��   Q���ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M���@Q�M�@x�ЋD�����E�P�I�I�ѡD��M�Q�@�@�Ѓ�Fu<�D���W�@�@`�Ћ�G�������3��D��EP�I�I�у���_^[��]Ëu��������������U���SVW�}����   �]���$    �D��ϋ��   �@��;���   =�m u~���( ����tq����� ��uV�E��E�    Ph�  ���E�    �v �D��M�Q���   �@X��SP�k������M����D�Q���   � uW�Ѓ���� ����u��D��ϋ��   �@4��SP�(�������u*�D��ϋ��   �@(�Ћ����%���_^3�[��]��Ѓ�_^�   [��]������������U��M��VW�@ ����ty�}��$    ��� ��uV�E��E�    Ph�  ���E�    � �D��M�Q���   �@X��WP�{������M����D�Q���   � u�Ѓ���� ����u�_3�^��]��Ѓ��   _^��]����������U��fnE��������} �YEt�E��E��$�] �]��,E�����]��E��E��$�d\ �]��,E�����]������U����M�V��� �E�Phacpihbyek�� �D��M���@j haqpi���   �Ћ��M�#u�� ��^��]��������������U���x  ����E�����E��E���   f.�����D{�M����^��   �E��U���   f.�����D{�E����^��   �E��M���   �U�E���E�}���   �M��$��L �} ��   �M�I �E؋U���   �������E���   �������M��*�������U��*B�������E�P�M�Q�U�R�M��L �*E��*M��^��\������^������E�\��   �YE��M��*E��*M��^��\������^������U�\��   �YE��E�@��	  �M��`Q�UR��X���P��Y  ����X����Y�X�����h����Y�h����X����$�_ ���]��E�f.�����DzH�M������`���f/��v�U����B��E����@�C  ��X����^EЃ��$�md  ��ݝ�����������^@��M����f/�h���v�U����\�E� �M�U��\��   �E� �M���   f/��v)�U���f/v�E� �X���M��<�U���f/��   v'�E� f/��v�M��\���U��E� �YE��M���`����^EЃ��$�c  ��ݝ�����������^(��U�B�E�@�\���M�X��   fW`��YE��U�B�  �E��`P�MQ��p���R�W  ����p����Y�p����M��YM��X����$��\ ���]��E�f.�����DzH�E���� ��x���f/��v�M����A��U����B�   ��p����^Eȃ��$�Ob  ��ݝ8�����8����^@��E� ���f/E�v�M����\�U���x����^Eȃ��$�0b  ��ݝ ����� ����^(�����\ȋE�H������Q�����R�E� �Y@����$�i[ ������Y������M�YA�X���U�\��   �YE��E� ����Y�����M�YA�X���U�\��   �YE��E�@�  �M��`Q�UR��@���P�U  ����@����Y�@�����P����Y�P����X����$��Z ���]��E�f.�����Dz�M�����  ��@����^E����$�`  ��ݝ�����������^@��U����f/�P���v�E����\ �M��U�E��\��   �M��U���   f/��v)�E���f/ v�M��X���U��<�E���f/��   v'�M�f/��v�U��\���E� �M��YE��U���H����Y���\���E�X��   fW`��YE��M�A��  �U��`R�EP������Q��S  ���������Y���X���U�\��   �YE��E� �������Y���\���M�X��   fW`��YE��U�B�o  �E��`P�MQ�U�R�{S  ���E��`P�MQ�U�R�tT  ���E��$�_  ��ݝ ����� ������M��$��������^  ��ݝ����������f/�����vj���E��$�^  ��ݝ�������������M��$��0����^  ��ݝ(�����0���f/�(���v	�E�    ��E�   �h���E��$�@^  ��ݝ�����������M��$������^  ��ݝ���������f/�����v	�E�   ��E�   �E�E�}� t�}���   �}��T  ��  ���f/E�v6�E�fW`��Y���X���M�\��   �YE��U��,�E��Y���X���E�\��   �YE��M��E��Y���\���U�X��   fW`��YE��E�@�J  ���f/E�v/�E��Y���X���M�\��   �YE��U�B�5�E�fW`��Y���X���E�\��   �YE��M�A�E��Y���X���U�\��   �YE��E� �   ���f/E�v.�E��Y���X���M�\��   �YE��U��4�E�fW`��Y���X���E�\��   �YE��M��E��Y���\���U�X��   fW`��YE��E�@�M���   ��t	�   �[�Y�E� f/��r>�M���f/r-�U�Bf/��r�E���f/@r	�E�   ��E�    �E���]ÍI nF +H �H A +H ]B �D �����������̡D���  � P���;��@����������U��D��M��� �@VW�u�@(Q�ЋD����}W�I�I�ыD�WV�A�@�СD��M�Q�@�@�СD����ϋ@�@<�Ћu;���   ���D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M��� �@�@<�ЋD�j�j�W�Q�M�P�BL�СD��M�WQ�@�@�СD��M�Q�@�@�СD��M�Q�@�@�ЋD����Q�ϋR<��;��6�����_^��]���������������U��D���0�@VW�}�@W�СD�j j�h���@W�@��j�E�h�  P�p����ȡD�WQ�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�@�E�jj
P�������M�D�Q�@�@�СD��M�Q�M�Q�@�@�СD��M����@�@<�ЋȡD�j��@�@Lj�VQ�M��СD��ϋ@�@<�ЋȍU�D�j�j�R�@Q�ϋ@L�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@��j�E�j
P�,������M�D�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���8�@�@<�ЋȡD�j�j�V�@Q�M��@L�СD��ϋ@�@<�ЋȍU�D�j�j�R�@Q�ϋ@L�СD��M�Q�@�@�СD��H�E�P�I�ыD��E�P�I�I�у���_^��]��U��D���0�@VW�}�@W�СD�j j�h���@W�@��j�E�jP�3����ȡD�WQ�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�@�E�jjP��������M�D�Q�@�@�СD��M�Q�M�Q�@�@�СD��M����@�@<�ЋȡD�j��@�@Lj�VQ�M��СD��ϋ@�@<�ЋȍU�D�j�j�R�@Q�ϋ@L�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@��j�E�jWP��������M�D�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���8�@�@<�ЋȡD�j�j�V�@Q�M��@L�СD��ϋ@�@<�ЋȍU�D�j�j�R�@Q�ϋ@L�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ��} ��   �D��M�Q�@�@�СD��M�j j�h���@Q�@�ЍE�P�O������M�D�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���$�@�@<�ЋȡD�j�j�V�@Q�M��@L�СD��ϋ@�@<�ЋȍU�D�j�j�R�@Q�ϋ@L�СD��M�Q�@�@�СD��H�E�P�I�ыD��E�P�I�I�у���_^��]�����U��D��M����@Q�@�СD��M�j j�h���@Q�@�ЍE�P�6^ �D��M�Q�@�@�Ѓ���]���������������U��D��M����@Q�@�СD��M�j j�hܲ�@Q�@�ЍE�P��] �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h��@Q�@�ЍE�P�] �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�L�E�P�I] �D��M�Q�@�@�Ѓ���]��U��D��M���`�@VQ�@�СD��M�j j�h$��@Q�@�СD��M�Q�@�@�СD��M�j j�h(��@Q�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��MЃ�4�@�@<�ЋD�j�j��Q�MQP�MЋBL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�ЍE�j P�����D����E�P�I�I�ыD��A�M�Q�M�Q�@�СD��M����@�@<�ЋD�j�j�V�Q�M�P�BL�ЍE�P��[ �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M��@�@Q�СD��M�Q�@�@�СD��M�j j�h0��@Q�@�ЍE�P�K����D����E�P�I�I�ыD��A�M�Q�M�Q�@�СD��MЃ�@�@�@<�ЋD�j�j�V�Q�M�P�BL�ЍE�P��Z �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ�^��]���U��D��M��� �@Q�@�СD��M�j j�h(��@Q�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M��� �@�@<�ЋD�j�j��Q�MQP�M��BL�ЍE�P��Y �D��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���]����������U���SV3�h�   Sh ��]���L h ��i� h�   h�  h �h�� 蠤 �� ��twjh�h�   j��A ������t���@ � ��3��D��M�Q�@�@�СD��M�j j�h`��@Q�@��V�E�   h    P�v �� ��t���3���t�D��E�P�I�I�у���^[��]���������������U��� j#h/� �@ ������   �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@��hƖ� j �E�P�E�Ph0� h/� �� �D��M���@�@Q�@�СD��M�Q�@�@�Ѓ��   ��]���������������U��E���   ����V��i�|  ��] �$��\ �E^�    �@   ��]ËE^�    �@   ��]ËE^�    �@   ��]ËE^�    �@�   ��]ËE^�    �@    ��]ËE^�    �@x   ��]ËE^�    �@   ��]ËE^�    �@
   ��]ËE^�    �@    ��]�(���EЋMfE�P����E��e6  �E^��]�(p���p����Mf�p���P����E��26  �E^��]�( ��E��MfE�PW��E��
6  �E^��]�(����@����Mf�@���P�����P�����5  �E^��]�(���E�MfE�P����E��5  �E^��]�(��E��MfE�P�P��E��z5  �E^��]�(@��E��MfE�P����E��M5  �E^��]�(����X����Mf�X���P�H���h����5  �E^��]�(����(����Mf�(���P�p���8�����4  �E^��]ËE^�     �@    ��]�IZ ^Z sZ �Z �Z �Z �Z �Z 3[ f[ �Z [ �[ �[ �[ \ K\ �\ �\   	
��������������U���\V�tY �D���h&� �A�ʋ@T�Ћ�����  �M��{d ���DY �D���Vh&� �A�ʋ@D�ЍM��d �Y �D���h&� �A�ʋ@T�Ћ���u^��]áD��M��E�   �E�   Q���   �@8�ЋD����Q��PhM  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��PhR  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��RhN  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����QP�B4��hO  �СD��M�Q���   � �СD��M��E�   �E��   Q���   �@8�ЋD����Q��PhP  �B4�СD��M�Q���   � �СD��M��E�   �E�    Q���   �@8�ЋD����Q��PhQ  �B4�СD��M�Q���   � �СD��M��E�   �E�x   Q���   �@8�ЋD����Q��PhS  �B4�СD��M�Q���   � �СD��M��E�   �E�   ���   �@8Q�ЋD�����ҋA��Rh]  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��PhT  �B4�СD��M�Q���   � �СD��M��E�   �E�
   Q���   �@8�ЋD����Q��PhU  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��Rh\  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��Ph_  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��RhZ  �΋@0�СD��M�Q���   � �СD��M��E�   �E�    Q���   �@8�ЋD�����ҋA��Rh[  �΋@0�СD��M�Q���   � �Ѓ�(���E�fE��M����P�E���.  �D��M�Q���   �@@�ЋD����Q��Ph^  �BH�СD��M�Q���   � ��(p��E����M�fE����P�E��.  �D��M�Q���   �@@�ЋD����Q��PhW  �BH�СD��M�Q���   � ��( ��E����M�fE�W�P�E��(.  �D��M�Q���   �@@�ЋD����Q��PhX  �BH�СD����   �M�Q� �СD��M��E�   �E�   Q���   �@8�Ѓ��M�fn��D����QhY  ��f�E��E��@�@H�СD��M�Q���   � ��(���E����M�fE����P�E��[-  �D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE����P�E���,  �D��M�Q���   �@@�ЋD����QP�BH��h�  �СD��M�Q���   � ��(��E����M�fE��P�P�E��,  �D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(@��E����M�fE����P�E��#,  �D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE��H�P�E��+  �D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE��p�P�E��S+  �D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � �Ѓ���^��]����������U�������u0�m(f(��]f(��e�\��}�\��M �\��\��Y��Y��$�Y��X�f(��Y��X�W��^�f/�w.f/��v�]�e �f(��Y$�Y��X��X�(��\��\��Y��Y��X�(��y4 �$�$��]��������������U��D�j �u�@@�@8�Ѓ�]�������U��M��t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ�]�3�]���������������^ ������    ������������h���^ �����    �=�� th����> �����    ���������U����D����VW���   �@X�Ћ��u�����   �}���D����   �΋@(�Ћ���tMj �u���j-�9; �D��M�Q�@�@�СD��M�j j�h\��@Q�@�СD��M�Q�@�@�Ѓ��D��M����   �@L�ЍE�P�a ���u����p���_^��]����������̡D����V3����   �@X�Ѕ�t�I �D�F���   �ȋR(�҅�u��^�����U��D����V���   �@X�Ѕ�t�u;�t�D����   �ȋB(�Ѕ�u�3�^]ø   ^]�������̡D����S���   �@X�Ћ؅�tzVW�3�W���6� ����t;�D����   ����RX�҅�t ��I ;�t#�D����   �ȋB(�Ѕ�u�j j W���� G��c|��D��ˋ��   �@(�Ћ؅�u�_^[��������U��=�� u3�]�VW�u������D����}3��ϋ��   ���   �Ѕ�~M��I �D���V���   ���   �ЋD�P���   ����Bh�СD���F���   ���   ��;�|������_�   ^]�����������U��=�� tuW�}��tl�D���V���   ���   �СD�������   �@X�Ћ���t9���$    ��D�V���   �ϋ��   �СD��΋��   �@(�Ћ���u�^_]��������������U��D��� �@VW���   �@��V�СD�j j�hP��@V�@�Ѓ��!� 3ɋ���D�VD��@�@�СD�j j�hT��@V�@�Ѓ��ۋ 3ɋ���D�VD��@�@�СD�j j�hX��@V�@�Ѓ��� 3ɋ���D�VD��@�@�СD�j j�h\��@V�@�Ѓ�菏 3Ʌ�D�jh��h�   j�E. ���� ��t���e, �|��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h`��@Q�@��V�E�Pj j �E�Ph� 莍 �D��M���@�@Q�@�СD��M�Q�@�@�СD�����@V�@�СD�j j�hh��@V�@�Ѓ��� 3ɋ���D�VD��@�@�СD�j �@�@j�hl�V�Ѓ��q� 3ɋ���D�VD��@�@�СD�j j�hp��@V�@�Ѓ��[� 3ɋ���D�VD��@�@�СD�j j�ht��@V�@�Ѓ��� j3Ʌ�h��h�   jD��, ���� ��t����* �|��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hx��@Q�@��V�E�Pj j �E�Ph� �� �D��M���@�@Q�@�СD��M�Q�@�@�СD�����@V�@�СD�j j�h���@V�@�Ѓ��]� j3Ʌ�h��h�   jD��+ ���� ��t����) �|��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@��V�E�Pj j �E�Ph� ��� �D��M���@�@Q�@�СD��M�Q�@�@�СD�����@V�@�СD�j j�h���@V�@�Ѓ��Ń 3ɋ���D�VD��@�@�СD�j �@�@j�h��V�Ѓ��� 3ɋ���D�VD��@�@�СD�j j�h���@V�@�Ѓ��9� j3Ʌ�h��h�   jD��O* ���� ��t���o( �|��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@��V�E�Pj j �E�Ph� 蘉 �D��M���@�@Q�@�СD��M�Q�@�@�СD�����@V�@�СD�j j�h���@V�@�Ѓ��a� 3ɋ���D�VD��@�@�СD�j �@�@j�h��V�Ѓ��;� 3ɋ���D�VD��@�@�СD�j j�h���@V�@�Ѓ��� 3ɋ���D�VD��@�@�СD�j j�h���@V�@�Ѓ��o� 3ɋ���D�VD��@�@�СD�j j�h���@V�@�Ѓ�虃 ��3Ʌ�D���_^��]��������VW艤 �����车 ���#��� ���#��g� ���#��ܱ ���#��� ���#�膸 ���#���� ���#��0� ���#��e� ���#��� ���#��� ���#��T� ���#��� ���#��� ���#��3� ���#��h� ���#��]� ���#��� ���#��W� ���#���� ���#��a� ���#��&� ���#���� ���#���� ���#��� ���#��� ���#��� ���#��Թ ���#��Y� ���#��N� ���#��3� ���#���� ���#���� ���#��b� ���#��G� ���#���� ���#���� ��_�#�^���������VW�y� ������]� ���#��B� ���#��'� ���#��� ���#���� ���#���� ���#��� ���#��� ���#��  ��_�#�^�������������U��U��u�A5 �Ѕ���   �D�h-� R�AL���   �ЋЃ���to�D�Vj R�A@�@8�Ћ�����tSW����  ����tDW���V�  ����t6S�]j ���� ��t�D���V���   ���   ��W����� ����u�[_^]�������U����D�VW���   ���   ���u�E�P�)����u��M�3���9}�   E��ޥ PWVh+� �� ���M��f� �D��M�Q���   ���   �Ѓ�_^��]�������U��E��dt8HtHu+�����t!Pj��o ]��Et�����tj��o �   ]Ë����t�D��q�@P�@�Ѓ���u�3�]���������Vjh��jej�$ ������t���o ����F    �5���
���    h�  hR� j h�u �= ���   ^�V�5����t �������n V��$ �����    hR� j �= ��^�����U��D�SV�u�@@�ً@,�ЋD������Q��j h�  �Rp�ҋD�j h�  �A�΋@4���u���,� ^�   []� �U��E��t	�E]�\U �D�V�u���   �N�@��-�� t��t��&t�F    3�^]� �F   �   ^]� �����U��W��� t.�O��t'�D�j Q�@@�@8�Ѓ��ȋj �u�w�RD_]� �D�SV�u�@@V�@,�ЋD����΋؋��   �RT�ҋD�j Ph�  �Q�ˋBl�Ћ���u�G^[3�_]� �D��΋��   �@��=�� u�w�   �D��΋��   �@��=�� �D�u!�@��j h�  ���   ���  P��  �6���   �΋@��=մ u0�D���h  h�  �@���   ��P�K�  ����P�p� �G�O���H����D�j Q�@@�@8�Ѓ��ȋj �u�w�RD^[_]� ���������V��N��t�D�j Q�@@�@8�Ѓ��ȋ�v�RL^� �����U��V��N��t-�D�j Q�@@�@8�Ѓ��ȋj �u�v�uV�RH��^]� �EW�^ �@]� ���U��Q�D�VW�}�@@W�M��@,�ЋD��������   �ϋRT�ҋD�j Ph�  �Q�΋Bl�ЋM��j �
� � -�  tL��t�u�M��u�u�uW�'S _^��]� ��tP�D��΋��   �@��3�=մ _����^��]� ��t&�D��΋��   �@��3�=�� _����^��]� _3�^��]� �U���E   V��t�U�B    �B    ��u��� �U�F�B�B   �u���u�u�uR�R ^]� �������������U��D��M�@�@ ��=neoa��   VW=ateg��   ��. �Ѕ���   �D�h-� R�AL���   �ЋЃ���t�D�j R�A@�@8�Ћ�����te����  ����tXW����  ����tJS�]j ���4� ��t�D���V���   ���   ��W���� ����uϋE[_^�    �@   ]ËE_^�    �@    ]ËE�    �@   ]��U���hS�]VWS�N� �D����E�P�I�I�ыD��A�M�QV�@�СD��M���@�@<�Ѕ��  �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�SQ�@�@(�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M̃�8�@�@<�ЋD�j�j��Q�M�QP�M̋BL�ЍE�P�k5 �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ�3��q  �}W��� �D����E�P�I�I�ыD��A�M�QV�@�СD��M܃��@�@<�Ѕ��D��@u~�@�M�Q�СD��M�j j�h���@Q�@�ЍE�WP�bC P�E�P�E�P�  P�4 �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ�83��  �u�΋@<�Ѕ���   j VS�F� ������   �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M�j j�h$��@Q�@�Ѓ�(�E�P�E�P�E�P�E�P�  ��P�E�P�  P�3 �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ� 3��  �D��M�Q�@�@�СD��M�j j�h8��@Q�@�Ѓ��E��M�P�RO j j �0�E��uj PS��N ���M������MP �D��M�Q�@�@�СD�����ti�@�M�Q�@�СD��M�j j�h$��@Q�@�ЍE�P�E�P�E�P�  P�2 �D��M�Q�@�@�СD��M�Q�@�@�Ѓ�,3��  �@���j h�~ ���   �ЋD����Q�M܋R<�҅���   ���E܋�P�F  �5�������Ѓ���t�D��A�M�Q���   �M��FB �D��M�Qj�M��@�@8�СD��M�Q���� V�@�M��@8�СD��M�Q���V�@�@8�СD�����P�EP���� P�B4�СD�����P�E�P���� P�BD�ЍM����B �U�D��M�Q����@�@8���� V�СD��M�Q���V�@�@8�СD�����P�EP���� P�B4��G���@�����d|0j hD��M��@  �E�P�1 �D��M�Q�@�@�Ѓ�3���D����Wh�~ �@�@4�о   �D��M�Q�@�@�Ѓ��D��E�P�I�I�у���_^[��]����������������U��D��M��4�@SQ�@�СD��M�j j�hX��@Q�@��j �E�Ph-� �N� ���M�D�Q�Ë@�@�СD��M��$�@Q�@�СD��M�j j��@�@��t,hh�Q�ЍE�P��/ �D��M�Q�@�@�Ѓ�3�[��]�h��Q��j j h�  h � j�E�Ph-� 蜑 ���M�D�Q�Ë@�@�СD��M��4�@Q�@�СD��M�j j��@�@��t,h��Q�ЍE�P�k/ �D��M�Q�@�@�Ѓ�3�[��]�h��Q��j j j h�� j �E�Ph*� ��J ���M�D�Q�Ë@�@�СD��M��4�@Q�@�СD��M�j j��@�@��t,h��Q�ЍE�P��. �D��M�Q�@�@�Ѓ�3�[��]�h��Q��j �E�Ph)� 詊 ���M�D�Q�Ë@�@�Ѓ�$��������D��M�Q�@�@�СD��M�j j�h���@Q�@�ЍE�Ph�� h�.  h�� �������M�D�Q�Ë@�@�Ѓ�(���;���j h���M��E  �E�Ph�� h�.  h�� �m������M�D�Q�Ë@�@�Ѓ��������j h��M���  �E�Ph � h�.  h�� �%������M�D�Q�Ë@�@�Ѓ��������j h��M��  �E�PhЪ h�.  h̴ ��������M�D�Q�Ë@�@�Ѓ����c���j h��M��m  �E�Ph � h�.  h�� �������M�D�Q�Ë@�@�Ѓ�������j h$��M��%  �E�Ph � h�.  h�� �M������M�D�Q�Ë@�@�Ѓ��������j h,��M���  �E�Ph�� h�.  hʴ �������M�D�Q�Ë@�@�Ѓ��������j h4��M��  �E�Ph�� h�.  h�� �������M�D�Q�Ë@�@�Ѓ����C���j h<��M��M  �E�Ph�� h�.  hѴ �u������M�D�Q�Ë@�@�Ѓ��������j hD��M��  �E�Ph0� h�.  h�� �-������M�D�Q�Ë@�@�Ѓ��������j hL��M��  �E�Ph@� h�.  h�� ��������M�D�Q�Ë@�@�Ѓ����k���j hT��M��u  �E�Ph�� h�.  h�� �������M�D�Q�Ë@�@�Ѓ����#���j h\��M��-  �E�Ph�� h�.  h�� �U������M�D�Q�Ë@�@�Ѓ��������j hh��M���
  �E�Ph�� h�.  h�� �������M�D�Q�Ë@�@�Ѓ��������j hp��M��
  �E�Ph� h�.  h�� ��������M�D�Q�Ë@�@�Ѓ����K���j h|��M��U
  �E�Ph�� h�.  h�� �}������M�D�Q�Ë@�@�Ѓ�������j h���M��
  �E�Ph� h�.  h�� �5������M�D�Q�Ë@�@�Ѓ��������j h���M���	  �E�Ph@� h�.  h�� ��������M�D�Q�Ë@�@�Ѓ����s���j h���M��}	  �E�Ph � h�.  hϴ �������M�D�Q�Ë@�@�Ѓ����+���j h���M��5	  �E�Ph�� h�.  h�� �]������M�D�Q�Ë@�@�Ѓ��������j h���M���  �E�Ph0� h�.  h�� �������M�D�Q�Ë@�@�Ѓ��������j h���M��  �E�Ph@� h�.  h�� ��������M�D�Q�Ë@�@�Ѓ����S���j h���M��]  �E�Ph� h�.  h�� �������M�D�Q�Ë@�@�Ѓ�������j h���M��  �E�Ph�� h�.  hմ �=������M�D�Q�Ë@�@�Ѓ��������j h���M���  �E�Ph`� h�.  hT� ��������M�D�Q�Ë@�@�Ѓ����{���j h���M��  �E�Php� h�.  hN� �������M�D�Q�Ë@�@�Ѓ����3���j h���M��=  �E�PhP� h�.  hִ �e������M�D�Q�Ë@�@�Ѓ��������j h��M���  �E�Ph0� h�.  hO� �������M�D�Q�Ë@�@�Ѓ��������j h��M��  �E�PhP� h�.  hʹ ��������M�D�Q�Ë@�@�Ѓ����[���j h��M��e  �E�Ph�� h�.  hش �������M�D�Q�Ë@�@�Ѓ�������j h ��M��  �E�Ph� h�.  h�� �E������M�D�Q�Ë@�@�Ѓ��������j h,��M���  �E�Php� h�.  hU� ��������M�D�Q�Ë@�@�Ѓ��������j h8��M��  �E�Ph�� h�.  h״ �������M�D�Q�Ë@�@�Ѓ����;���j hD��M��E  �E�PhP� h�.  hQ� �m������M�D�Q�Ë@�@�Ѓ��������j hL��M���  �E�Ph � h�.  hԴ �%������M�D�Q�Ë@�@�Ѓ��������j hX��M��  �E�Php� h�.  hд ��������M�D�Q�Ë@�@�Ѓ����c���j h`��M��m  �E�Ph� h�.  hP� �������M�D�Q�Ë@�@�Ѓ�������Vjhh�h�   h�  �} ����t���O  ���3�j h@��M���  j h8��M���  j h���M���  �E�P�M���? V�M�Q�0�E�j Ph&� ��k ���M������@ �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���tj h���  jhh�h�   j � ����t���B  ���3�j h���M��-  j h8��M��  j h���M��  �E�P�M���> V�M�Q�0�E�j Ph�� �k ���M�������? �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���tj h����   jhh�h�   j��
 ������t���	 �|��3�j h���M��Z  j h��M��K  V�E�Pj j �E�Ph� �dj �D��M�Q�@�@�СD��M�Q�@�@�Ѓ� �M�j h��   h�z �E�Ph+� �-� ���M̡D�Q�Ë@�@�Ѓ�j ��t2h��M���  �E�P�! �D��M�Q�@�@�Ѓ�^3�[��]�h8��M��  j hH��M��  j j �E�Ph� j �E�Ph.� �� ���M̡D�Q�Ë@�@�СD��M�Q�@�@�Ѓ�$��u�j hX��M��&  j h���M��  hƖ� h/� �E�P�E�Ph � h'� �6� ���M̡D�Q�Ë@�@�СD��M�Q�@�@�Ѓ� 3�����^[��]����������������U��V�u��V�    �F    �D����   �@�Ѓ���^]� ���������������U��V�u��V�    �F    �D����   �@$�Ѓ���^]� ���������������U��D�V��V�@�@�СD�V�u�@�@�Ѓ���^]� �U��D�V��V�@�@�СD��uj��@�uV�@�Ѓ���^]� ������������U����   V���?V h����<����H��F    �F    ��
 Ph����t����
 Ph���M��
 P�E�P��, ��P�E�P�5 ��P��X���P�% ��P�E�P� ����X����* �M��" �M�� �M�� ��t���� ��<�����
 �=�� u��D j j��M���Q���zA �M���
 ��^��]������������V���H �N�T��
   ��^�������U��QSVW���2e �K���������KD�����Kx�����ˍ��   �G   �C�Kj jh���P8�CD�KDj jh ��P8�Cx�Kxj jh���P8_^��[��]���������VW���T ����w ���W�NN�F(O`Op��   ��   ��   ��   ��   Ǉ�      Ǉ�       Ǉ�   ����Ǉ�       Ǉ�       Ǉ�      Ǉ�       Ǉ�   ����Ǉ�       Ǉ�       Ǉ       Ǉ      Ǉ      Ǉ      Ǉ  ����Ǉ  �����  �(  �h����F�>�^����G�ǉw�_^�U���SVW��� ���s�D�V�@�@�СD��{ W�@�@���1 �C�M�D�Q�@�@�СD��M�j j�hx��@Q�@�СD��M�VQ�@�@�СD��M�Q�@�@���0 �C�M�D�Q�@�@�СD��M�j j�h���@Q�@�СD��M�WQ�@�@�СD��M���D�@Q�@�Ѓ�_^��[��]��������������V���ȵ �����F8W�����F@�FH   �FL�F\�Fl�F|���   ���   ǆ�       ^�����V���h� ( �W��p����<�V`Vp��   ��   �F4    FP�F8   W��F<    �F`ǆ�      (0��FxW�f�Vp���   V@f֎�   f֖�   ^������������VW��� �O����a �O�G|��h ��_^�����̡D�V��V���   ���   �Ѓ��    ^���������������V�񍎰   W�������5Q j �Nx�FxH��U �=�� th���a@ ���Nx�Q j �ND�FDH��uU �=�� th���2@ ���ND��P j �N�FH��FU �=�� th���@ ���N�P _��^�` ����������������� �����������U���   �M�y8�iXf(��A@�YAP�q(�Q �Y��E�f(��M��\�f(��A�YIP�E�(��YQ@�Y��M�(��U��Q0�\��E�(��]��qH�Y��Y���x����M��\��E�(��Y�W��u��e��X�(��Y��X�f.џ��Dza�EW�HH H0H@HP� (���@(���@0f�HW�f�H(f�H@����@Hf�HX��]�����^��q�E�(��Y�(��YA@�if(��	�Y�(��YQP�E�f(��Yq(�\��Yi (��\��\��e��Y}��YA0�Y��X��E��\E��Y��X��E��\E��Y}��Y��}�(��\��\��o�x����Y}��X��oE��\��X��U��\U��o]��Y��Y}�f(��Y��I0�Y��X��Ya@�X��m��Y��Y���x����u��E��E�(��Y��YQX�E��E��Y��E�(��YAX�\�f(��YA(���YY(�Y��\��Y��YIP(ƋE�YA@f��\��E��YA8�Y��\��oE��YA �Y��E�f(�f��YAP�ou��\��u��oE��q0�Yq �Y��E��E��YA8�\��o�x����Y��m��E��oE��M�f�� �oE�f��@�E�f��oE��p �`0f��X@�@P��]���������������U��M�U�;u$�A;Bu�A;Bu�A;Bu�A;Bu3�]ø   ]�������U��M�E�I��`�A0�X�YʋE�Y��X	�X��AH�Y��X��A8�Y���I �Y��XI�X��AP�Y��X��A@�Y��H�I(�Y��XI�X��AX�Y��X��H]����������������U��D�V�uV�@�@�СD�V�u�@�@�СD����΋@�@<�ЋD�j�j��u�Q��P�RL�ҋ�^]������������U��M�E�I�`��A0�X�E�Y��Y��X��AH�Y��X��A8�Y���I �Y��X��AP�Y��X��A@�Y��H�I(�Y��X��AX�Y��X��H]��������������U��V��j �H��mO �=�� th���*: ������J �Et	V�� ����^]� ����������U��V���x��?� �Et	V��� ����^]� ���������U��V���P��� �Et	V�� ����^]� ���������U��V������߭ �Et	V�� ����^]� ���������U��V���ع语 �Et	V�S� ����^]� ���������U��V��N<�\���t踏 �F<    ���j� �Et	V�� ����^]� ����U��V���H��?� �Et	V��� ����^]� ���������U��V������� �Et	V�� ����^]� ���������U��V������߬ �Et	V�� ����^]� ���������U��V���h�诬 �Et	V�S� ����^]� ���������U��V������� �Et	V�#� ����^]� ���������U��V���0��O� �Et	V��� ����^]� ���������U��V������� �Et	V��� ����^]� ���������U��V������� �Et	V�� ����^]� ���������U��V�����迫 �Et	V�c� ����^]� ���������U��V��N��������� �Et	V�/� ����^]� �����U��V���u����Et	V�	� ����^]� ���������������U��V������G �Et	V��� ����^]� ���������U��V���p���� �Et	V�� ����^]� ���������U��V�����Ϫ �Et	V�s� ����^]� ���������U��V��F��P�$ �FP�$ �D��H�F P�A�СD��H�FP�A�Ѓ����� �Et	V�
� ����^]� U��V������?� �Et	V��� ����^]� ���������U��V���ؾ�� �Et	V�� ����^]� ���������U��V������ߩ �Et	V�� ����^]� ���������U��V����诩 �Et	V�S� ����^]� ���������U��V������� �Et	V�#� ����^]� ���������U��V�����O� �Et	V��� ����^]� ���������U��V���8��� �Et	V��� ����^]� ���������U��V������� �Et	V�� ����^]� ���������U��V����迨 �Et	V�c� ����^]� ���������U��V���T�菨 �Et	V�3� ����^]� ���������U��V���P��_� �Et	V�� ����^]� ���������U��V���<��/� �Et	V��� ����^]� ���������U��V�������� �Et	V�� ����^]� ���������U��V���%� �Et	V�y� ����^]� ���������������U��V�����蟧 �Et	V�C� ����^]� ���������U��V���H��o� �Et	V�� ����^]� ���������U��V���L��?� �Et	V��� ����^]� ���������U��V���,��� �Et	V�� ����^]� ���������U��V��N4�,���t�D��@ �@T���F4    ���¦ �Et	V�f� ����^]� ������������U��V���l�菦 �Et	V�3� ����^]� ���������U��V���<��_� �Et	V�� ����^]� ���������U��V������� �Et	V��� ����^]� ���������U��V�������� �Et	V�� ����^]� ���������U��V��N �� ���� �Et	V�o� ����^]� �����U��VW���O�G|��jY �O�R ����� �Et	W�/� ����_^]� ����U��V��N�|��,Y ����Q �Et	V��� ����^]� ���������������U��V�������= �Et	V��� ����^]� ���������U���Mf/��r��]����f/�r�(�]�(���� �E�E]���U����E� � �E��E���]�����U����EfTP��E��E���]��U���SVW��� �Ѕ�t7�D�h-� R�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3��D��M�Q�@�@�СD��M�j j�h$��@Q�@�ЍE�P�}
 ����t~�D�j����@V�@�СD��M�VQ�@�@�Ѓ����5� �ˋ��<D ���+�����P�D ���+�����P�.� ��������$��� V���?� �   �3��D��E�P�I�I�у���_^[��]���������Vjh��h6  j@�L� ������t%��謢 ������x��F4   �F8^�3�^�����������Vjh��h�  j`��� ������tE���\� (����F8�P�����FH   �FL    �FP�FX   �F\   ^�3�^�����������Vjh��h�   jx�� ������tY���� W����N8��NHNX�Fh   W��Fl   �F8( �f�NH����FPf�N`�Np^�3�^�������Vjh��jbjP�� ������t%���o� W��عN8��W��F8f�NH^�3�^��������������Vjh��h
  j@�� ������t&���� �\����F4   �F8    �F<    ^�3�^����������Vjh��h�  j<�l� ������t���̠ �H����F4    �F8    ^�3�^�Vjh�h2  jP�,� ������t5��茠 W�����F4    ���F8   �F@�FH   �FL    ^�3�^�����������Vjh��h�   jL��� ������t;���,� ������F4   �F8   �F<   �F@    �FD   �FH   ^�3�^�����Vjh��hc  j@�l� ������t%���̟ ������h��F4    �F8^�3�^�����������Vjh�h�  j`�� ������t@���|� (���F8���W��FP   �FH�FT   �FX   �F\    ^�3�^����������������Vjh��h  j`�� ������tA���� �����F8W��F@����0��FH    �FP�FX   ^�3�^���������������Vjh�h�  jH�<� ������t,��蜞 ���������F8�F@   �FD    ^�3�^����Vjh��h�   jh��� ������t'���L� W����F8��( �FHFX^�3�^���������Vjh��h�  jH�� ������t%����� ��������F8�F@    ^�3�^�����������Vjh��hQ  jX�L� ������t+��謝 (����F8�p�W��FP   �FH^�3�^�����Vjh��hR  h�   ��� ������tI���Y� W���F8���FP    �FHFX�Fx    �Fh����Fp���   ^�3�^����jh�h�  j0�� ����t������3��������������Vjh�h;  jH�\� ������t%��輜 � �������F8�F@   ^�3�^�����������Vjh��h�  h�   �	� ������tS���i� ( �W��ؾ���F4    �F8   �F<    �F@�NH�FPNX�FhNp��   ^�3�^����������Vjh��h�  jH�� ������t,���� � �������F8�F@    �FD   ^�3�^����Vjh�j`jX�?� ������t;��蟛 W����F@������F4    �F8    �FH�FP   ^�3�^��������Vjh��h�  j4��� ������t���<� �����^�3�^���������������Vjh��hs  j4�� ������t����� ����^�3�^���������������Vjh��jj@�_� ������t%��迚 ������8��F4    �F8^�3�^��������������jh��h�  h�   �
� ����t������3�����������Vjh�hB  j4��� ������t���<� ����^�3�^���������������Vjh�h�  jP�� ������t#����� ( ����T�F8�FH    ^�3�^�������������Vjh��jj4�O� ������t��诙 �P���^�3�^��jh�h  h�   �� ����t������3�����������Vjh�h�  jX��� ������tB���L� W�����F8������F4    �F@�FH   �FL   �FP    ^�3�^��������������Vjh��j.j�� ������t���� �����F    �F    ^�3�^����Vjh�h(  jP�<� ������t:��蜘 ���������F8�F@   �FD   �FH   �FL    ^�3�^������Vjh��jj@��� ������t&���?� �H����F4    �F8   �F<   ^�3�^�������������Vjh�h  j`�� ������t@���� (����F8�L�W��FP   �FH�FT   �FX   �F\    ^�3�^����������������Vjh�h%  j8�� ������t���|� �,����F4    ^�3�^��������Vjh��jj8��� ������t���?� �,����F4    ^�3�^�����������Vjh�h�  j4�� ������t����� �l���^�3�^���������������Vjh��jh�   �\� ������t7��輖 W��<�F8��FH�FX( �F`(`�Fp^�3�^���������VjhԵjaj��� ������t���� �����^�3�^��VjhT�h�  j4��� ������t���,� �����^�3�^���������������VjhT�jXj�� ������t���?� ����^�3�^��Vjh��jj�_� ������t���� �p���^�3�^��U��VWjh�jujH���)� ������t:���) �u��PV� V�O ����� W��G@    �G8�G_^]� _3�^]� ��������������U��D����   ���   ]�����������U���V���q �D��M�Q�@�@�СD��M�j j�h��@Q�@�Ѓ��E���P�q �D��M�Q�@�@�Ѓ���h�� ��q ���Rr h�� ����q h�� ����q h�� ���q h�� ���q ���r hô ���q ���r h�� ���q h�� ���q ����q h�� ���mq ���6q �D��M�Q�@�@�СD��M�j j�h$��@Q�@�Ѓ��E���P��p �D��M�Q�@�@�Ѓ���h�� �q ���vq hƴ ����p hĴ ����p hŴ ����p ���Kq hǴ ����p hɴ ����p ���,q h�� ���p ���yp �D��M�Q�@�@�СD��M�j j�h,��@Q�@�Ѓ��E���P�p �D��M�Q�@�@��h�.  ��K ����P��o hd� ���>p he� ���2p h�� ���&p ����o h�.  �K ����P�o hf� ����o hy� ����o hg� ����o hh� ����o hi� ����o hj� ����o h}� ���o hk� ���o ���so h�.  �9K ����P�.o hl� ���o hm� ���vo hn� ���jo ���3o h�.  ��J ����P��n ho� ���Bo hp� ���6o hq� ���*o hr� ���o hs� ���o h{� ���o ht� ����n hv� ����n ���n h�.  �}J ����P�rn hw� ����n hx� ���n h� ���n ���wn h�.  �=J ����P�2n h�� ���n h�� ���zn h�� ���nn h�� ���bn hz� ���Vn h�� ���Jn hu� ���>n h�� ���2n h�� ���&n h�� ���n h~� ���n h|� ���n h�� ����m ���m ���m �D��M�Q�@�@�СD�j j��@�@�M�h4�Q�Ѓ��E���P�Om �D��M�Q�@�@�Ѓ���h&� �m h'� ���m h(� ���wm h)� ���km h*� ���_m h+� ���Sm h,� ���Gm h-� ���;m h.� ���/m h/� ���#m ����l ���m ^��]�U���V���rl �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���P�il �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �l �D��M�Q�@�@�Ѓ�����l �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �Ql �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �l �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �k �D��M�Q�@�@�Ѓ����8k �D��M�Q�@�@�СD��M�j j�h��@Q�@�Ѓ��E�P����j �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �k �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  ��j �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E�Ph�  ���rj �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �#j �D��M�Q�@�@�Ѓ����Hj �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  ��i �D��M�Q�@�@�Ѓ�����i �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���Ph�  �qi �D��M�Q�@�@�Ѓ�����h ���i ^��]�����������U���W���? ��   SV�G�����G�, ����, �M�_W���Gfn�fn��������G�O ��tI�,�P�,�P�u� �M�wVS�ȶ �M蠷 ��]��M��Y��O(���Y��^[_��]� ��U��E��wT�$�D� ��  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]Ã��]��� ��  � � � ?� � � ?� #� ?� *� 1� 8� ����U��E��wQ�$��� 3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø
   ]Ã��]ÍI �� �� �� �� �� �� �� �� �� �� �� �� �� �� ����U��E��wT�$��� �@  ]øB  ]øC  ]øD  ]øE  ]øF  ]øG  ]øH  ]øI  ]øA  ]øL  ]Ã��]�2� 9� @� G� N� � U� \� � c� � j� q� x� ����U������  �EV��W�t$�    �~P �@    �@�����@    �@    �W  �� �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��vP�����  �D����NTj h\  �R�|$���   �ҋD��NTjhY  �R�D$d���   �҉D$X����  ��I �D�j W�@@�@8�Ѓ����t$;}�y  �|$\ ��   �L$��$�   WP�I ���  ��$�   ��$�   �Y����P�D$$��$�   �Y���D$<�q� �L$��$�   ��$�   � �X�\d$ �\\$8�AH�i(�Y��Y��Y��Y��A8�X�f/���  �X�f/���  �Q0�A@�X�f/���  �X�f/���  ���3��@d�Ѕ��y  �����W�@\�Ѕ��S  �L$W�� �D$,���=  �t$��$   W�t$�� P����  jc�t$0���o ��$  P�D$|�D$D��  �ЋD$X�T$0�o�D$H���c  �D$p�2   �\D$HW���$�   ��$�   ��$�   fTP��Y����$�   ��$�   ��$�   �,���2��Xl$PLȃ������l$Pfn��������$�   ��$�   ��$�   �D$(�L$(fn��������o�$�   ��$�   ��$�   �X���$�   �(��Xt$`f��X��L$(W��D$���o�t$H� �ă�����$�   f�� �ă���f�� �����$�   P�� �D$ �   ��$�   �D$8��$�   �D$�o�$�   ��$�   �D$H��$�   E�o�$�   D$`���$    �fnƃ�����L$H���^`��D$���o�L$@� �ă��o�$�   �I ��ă����� ��$�   P�Q� ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��l$�D$��$�   �f(��D$�D$`��\��T$h�\���\�f(��\�(��Y��Y��Y��X�f(��Y��X�W��^�f/�w)f/��v�l$f(��(��Y��Y��X��X��L$h�D$`�\��\��Y��Y��X��]� �H�f/���  �o�$�   F�o�$�   �o�$�   ��$�   ���]����y  ���q  �D$H�}�L$L�\$P�D$0�D$8�T$@�e�u�D$�D$<�|$p�|$0��m���L$8�L$��D$8�\��\$ �\$T�T$H�T$D��D$8�D$ �d$8��\$H�f(��D$ �\��\��|$0�|$p��L$�Y��D$Hf(��l$H�\�f(��Y��Y��X�f(��Y��X�W��^�f/�v�D$�-f/��v�D$0�\$ �(��Y��Y��X��XD$�\��\��Y��Y��X�f(��� �H�f/�wA�t$���G�@d��;�������|$�D$���pP臂 ���|$���I����E_^��]� �M�D$�A�D$,�y_�A���   ^��]� ����������U��D�S�]V�@@WS�@,�ЋD������Q��j h�  ���   �ҋD������   �ˋR��=�� ��   ����   �D���V�u�@h�  �@l�ЋЅ�tn�D�jR�AH���  �ЋD����؋Q��Vh�  ���   ��;�t8�D���Sh�  �@�@4�СD��MVhȴ ���   �@��_�F^[]� _��^[]� �������������U������   �ES��VW�\$�{P �    �@    �@�����@    �@    �o  ��� �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��sP����  �D����KTj hU  �R�t$���   �ҋKTj h\  fn��D�����@���   �D$x�Ћ��|$����  �D�j V�@@�@8�Ѓ���;u��  ����   �|$��$�   VP�O �.�  ��$�   ��$�   �Y����P�D$4��$�   �Y���D$衂 �GH��$�   ��$�   � �X�\d$0�\\$�o(�Y��Y��Y��Y��G8�X�f/���  �X�f/���  �W0�G@�X�f/���  �X�f/���  ���3��Pd����  ���W�P\���x  W���P� �D$D���d  �t$jcP��$�   P�N ��  W�t$�N �o ��$�   P�D$l��$�   �Ź  �]�}�u�o�e�T$P�l$P(��D$X��U����T$0��$�   �l$H�l$x�D$�T$ �T$H��l$(�ol$`�L$((��T$H��U�l$l��D$�\����L$(�T$`�oT$0�\$`�f(��D$0�D$�D$ ��l$0�\��\��D$ f(��\��Y�f(��Y��Y��l$0�X�f(��Y��X�W��^�f/�v�l$(�D$ �=f/��v�l$H�D$�%f(��YT$0�Y��XD$((��D$ �X�f(��\��\��Y��Y��X�f(��M� �L$pf/���   �L$P�D$X�\�$�   �\L$x�Y��Y��X��� �Y���L$P�\M�D$`�D$X�\E�Y��Y��X���� �\$pf(��D$`f(��X�f/�v
�\�f/�w@�t$���G�Pd;��h����|$�D$���pP�| ���t$���7����E_^[��]� �M�D$�y_�A�D$@^�A���   [��]� ���������������U���SV��W�FH�E�ǆ�      ǆ�   ������� �ȅ�t7�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3ۡD�j ���   �@@�@8�Ѓ����~P ��   ���    ��   ����PT����   ����Pd����   ���j �P\����   ���   j �| ����   P�E���P���   �L� ��ur�M�f�f.�����DzW����   f^�E�fE����   �΃���� �E�P������}�u"�oE�E����   ���   �   _^[��]�_^3�[��]��������������U���DSW�}3ۉ]�����  �D�h-� W�@L���   �ЋЃ�����  �D�SR�A@�@8�Ѓ��E����v  V�u��u���Hw  �����  9]��   �D��M�Q�@�@�СD��M�j j�hp��@Q�@�СD��M�Q�@�@�СD��M�j j�hD��@Q�@�Ѓ�(�E܋λ   j$P�Z� P�E�P�E�P�������P�E�P�������P�� ���E��t�E ��t�D��M�Q����@�@�Ѓ���t�D��M�Q����@�@�Ѓ���t�D��M�Q����@�@�Ѓ���t�D��M�Q�@�@�Ѓ��} t^_3�[��]� �M�WV�+  j j h�� ��� j j h,� ��� ���   ^_[��]� _3�[��]� �������VW���� �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��wP�����  ����tj���� �wP���x ����u�_^���������������U���,�}�  V����   �u�M���� ����' �D�Phdiem�Q�M�B4�СD��M�havem�@�@X�Ћ�M�Q���P@�D���Phavem�Q�M싂�   �СD��M�Q���   � �Ѓ��E��P�3' �M��� �   ^��]� ���������������U��E��|SVW��=�  ��   tl=�  �l  �D��u��j havem�@���   �Ѓ�d�G  �D���j j�@���   ��j P���5�  Ph�� ��� ���   _^[��]� j h�� �-� ���   _^[��]� F�������  �$��� ��� ����  jj P������_^�   [��]� �M��H� j hh��M��)���j hp��M������E�P�E�Pj j �M��V� ���MԡD�Q�Ë@�@�СD��M�Q�@�@�Ѓ���u7j �E�jP��� ���E��t �� ��tP�u���}�  �EP�� ���M��� _^�   [��]� ��� ����  �������  PQ���7�  _^�   [��]� �� ��V茐�������r  �E����  �M��?� j hh��M�� ���j hx��M������E�P�E�Pjj �M��M� ���M��D�Q�Ë@�@�СD��M�Q�@�@�Ѓ����*����f� �E��t&�u��PV��  ��thBF j�E�P�u�<� ���EP�@� ���E    �M��~� _^�   [��]� ��� ��V裏��������q  �؅���  �=�� th����� �����    ��� SPV�ϣ���K  _^�   [��]� �h� ��V�@��������fq  �؅��^  �=�� th���� �����    �g� SPV�ϣ����  j SV���m���_^�   [��]� ��� P�E�ю����������� ����  �M��� j hh��M��f���j hx��M��W����E�P�E�Pjj �M��� ���M��D�Q�Ë@�@�СD��M�Q�@�@�Ѓ����p����� �E���h������*�  ����t�]�V�u��S�  ��轝 ����u�hBF j�E�P�u�d� �EP�k� ���E    �M��� _^�   [��]� ��� ��S�΍����������� ����   �=�� th���� �����    ��� �Σ���y�  ������   V�5����S�`  ���	� ����u�_�F^[��]� �r� P�L��������ro  ����tn����� P�M�輷���E�P�� ����t:�E���P�A� j Vh�� �� �D��M�Q�@�@�Ѓ��   _^[��]� �D��M�Q�@�@�Ѓ�_^�   [��]�  � �� �� 3� �� �� �� �� )� ������������U���VW�� �����z� �D��E�P�I�I�ѡD��M�j j�h0��@Q�@�СD��M�Q�@�@�Ѓ��σ}cj uT�uVj*�e� �D��M�Q�@�@�СD��M�j j�h<��@Q�@�СD��M�Q�@�@�Ѓ�j�u�u�R�uVj*�� �D��M�Q�@�@�СD��M�j j�hH��@Q�@�СD��M�Q�@�@�Ѓ�j�u�u���v ���� �D��M�Q�@�@�СD��M�j j�hT��@Q�@�СD��M�Q�@�@�Ѓ�_^��]� �����U����oEVj �������(  � �E�P� �}�ue�M��E�9�  u9�  tm��  ��  9�  t��  cu��cu3���  ^��]� ��cu���=�  ���@��  ^��]� ǆ      ǆ  ����ǆ      ^��]� ����������������������U���$SV�uW�}��tRV�� �Ѓ����tB�D�RW�AT�@�Ѓ���t+����s �Ѕ�t�D����   �ʋ@��=.� ��  �]$��t8�D�h-� S�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E��E    �M��p �D�W�E�I@�I,��V�E�� h.� �E��Ur �����ˉu�j Vj,�� �D��A�M�Q�@�СD��M�j j�hx��@Q�@�СD��M�Q�@�@�Ѓ�����  �D�V�@@�@,�ЋD������Q���uh�  �Rp���u� �D�����0����A��Rh�  �@4��j Wj(���� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD����ϋ��   j �u����   �СD��u�W�@T�@�Ѓ����7r �E�����   �D����   �ȋRx�҃����D���W�S�@j�u���@����V�СD�VW�@�@�ЋM��h�� �#� ���D�W�@@�@,���oE����������t �D��]����   �ˋ@L��jW�u������M��P�r �D���j S���   ���   �СD���Sh�  �@�@p�СD��u��u��p������M��P�Fp��_^[��]�������������U���l�D�SVW�@@�u�@,�ЋD��u�E�I@�I,�ыu$��3��E�}���I W� ��S�$  �D����E�Q�M�j S���   �҅��  �E9E��  j �E��E�    PS�M��E�    ��: �MP�� �M���< h.� V�M��Ŷ ����  ��t8�D�h-� V�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E���E�    �M�m h.� �E���n ���E��j Pj,�S� �D��A�M�Q�@�СD��M�j j�h ��@Q�@�СD��M�Q�@�@�ЋM���D����"  �@@Q�@,�ЋD������Q���uh�  �Rp�ҋD�Sh�  �A�΋@4�Ћu$��j �uj(�� �D��M�Q�@�@�СD��M�j j�h,��@Q�@�СD��M�Q�@�@�СD����M���   j �u��   ��j �E��E�    PS�M��E�    �/9 �MP�v� �M��.; hK  V�M�� � �E�����   �D����   �ȋRx�҃����D���W�V�@j�u���@����V�СD�VW�@�@�ЋM���h�� �� ���D�W�@@�@,���oE����������Eq �D����   �M��@L��jWS�x  �M��P�<o �D���j �u����   ���   �СD����u�h�  �@�@p�Ћu$�}�D��u�M�S�@�@p�СD��M�Q���   � �Ѓ��D��M�Q���   � �Ѓ�G�}���H�����_^[��]Ë��   �M�Q� �Ѓ�_^[��]����������U���SV��W�]��� ����t7�D�h-� W�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3��y� �E��D����   ���   �ЉE��E����  �D�WP�I|�A$�Ѓ�����   �sP��� y  �]������   �I j ���i ��t�D����u�j ���   � �Ћ���tLj Wj,���۾ �D��A�M�Q�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��D��M�W���   ���   �ЋE���pP�h �����]����D��M����   ���   �Ѕ�tjS�u�躄���D�j�u��@|�@,�Ѓ��J�D��M�Q�@�@�СD��M�j j�h`��@Q�@�ЍE�j P�]� �D��M�Q�@�@�Ѓ� �D��M�Q���   ���   �ЍE��E�    P��� ��_^[��]� ������U��Q�D�V�u�u���   �u�M��v�I�@�СD��u�M��u���   �v�I�@�и   ^��]� ��������������U���S�]W���.  �D�h-� S�@L���   �ЋЃ����  �D�j R�A@�@8�Ћ�������  �U����  �D�h-� R�AL���   �ЋЃ�����  �D�j R�A@�@8�Ѓ��E�����  V�� �E���u  �D�SP�I|�A$�Ѓ����Z  �D��u�u��j ���   � �ЋM�jP�E��� V���u  ������   ���$    �D��uj ���   �ϋ ���u�ȉE��,l �D��E��u����   �H�Rh�ҡD��ϋ��   �@��-�� t��&uy�D�W�@@�@,�Ѓ���Sh�  �F� �Ѕ�tU�D��uj ���   �ʋ �ЋM��j j V�
� �D��u��I@�I,�ыD����ЋA��Vh�  �@p�ЋuV���sd ���������D�j�u�@|�@,�Ѓ��E�   P�V� ����^_[��]� �E3�P�=� ����^_[��]� _3�[��]� �����U��E=Ҵ u	�E]� �E���   ]�;   ����������̸   � ��������U��}�� u�O�  �   ]� ������U���@SVW���p� �u����w� �  ��d� �7  ���� ��   tD��,� �  ���� �  ���� �  �{P �  V���ϐ �   _^[��]� �{P ��  �D��Mj h1icM�@���   �ЋD����Mj h2icM�R���   ��j PWh���h������{� �   _^[��]� ��CK�����z  ���� �$��� h���h�������� �   _^[��]� ���ʽ���   _^[��]� ��� �T  �r  ��x� ��   �  ��~� �  ����� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��E���jP�ia  �����o V�����  P���<  ��襸 �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��   _^[��]� hG  ���  ���0  ���� ����j hl��̦���WQ�����E���jP�`  �����o hx� ����>  P���
  ���� ����j hx��~����	Q�����   _^[��]� h�� ���,  ����  ��荷 �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��EЋ�jP�`  �����o h� ����  P����	  ���9� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��   _^[��]� ��cdpu��   ��   ���C������   ���� �$��� W�z��������   ���\  ����   9CP��   P���<� �   _^[��]� �D��Mj h1icM�@���   ��P���� �   _^[��]� jW覇��W� z������t%���B\  ��t9CPtP�j ���ͥ j ���t� _^�   [��]� ��� ?�  � �� ��          ��� �� "� ��           ���U��E�C����(�]  �$�X� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� �ʴ ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� ��� ]� �̴ ]� �ʹ ]� �ϴ ]� �д ]� �Ѵ ]� �Դ ]� �մ ]� �ִ ]� �״ ]� �ش ]� �N� ]� �O� ]� �P� ]� �Q� ]� �T� ]� �U� ]� �S� ]� ���]� �� � � � � (� 1� :� C� L� U� ^� g� p� y� �� �� �� �� �� �� �� �� �� �� �� �� �� �� Q� Q� Q�  � 	� � � $� -� 6� ?� H� ����U���SVW���0	 �D��؍E�P�R�R�ҋD�j j�h@��A�M�Q�@�Ѓ��E���P� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���j j j Pj jj?h�  �2 �D��M�Q�@�@�Ѓ���j �+3 jjjj���L3 jj���2 �E�����j j j?h�  ���h0 �E����   j �E���PV�0 ���Z2 ���1 jjj h�  ���E������*0 �E���j �E�P�GP�f0 �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���j Pj jjj �( �D��M�Q�@�@�Ѓ��E�������jjj h�  �/ �E���j �E�P�GDP��/ �D��@�@�M�Q�СD��M�j j�h���@Q�@�Ѓ��E���j Pj jjj �' �D��M�Q�@�@�Ѓ��E�������jjj h�  �"/ �E���j �E�P�GxP�^/ �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���j Pj jjj �' �D��M�Q�@�@�Ѓ�����0 ����P$����P_^��[��]����������j jxj h�  �`( �   �����������U���VW���A �D����E�P�R�R�ҋD�j j�h���A�M�Q�@�Ѓ��E���P�	 �D��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E���j j j Pj jj?h�  �/ �D��M�Q�@�@�Ѓ���j �<0 jjjj���]0 jj����/ j j j?h�  ���+ h�  W�O� ���{/ ���4���_��^��]�������������U���$SVW��耵 �D��KTjhZ  �R�E����   �҅���  �uV�a� ��������  �D������� ��@V�@tD�СD�j j�h���@V�@�Ћu��E����VP耗  �D�P���   �ϋB|�ЍM��B�СD�j j�h���@V�@�Ћu��E܃���VP�<�  �D�P���   �ϋB|�ЍMܡD�Q�@�@�Ѓ����m� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ���j j W�ҙ j Wj,���V� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@��j �� ����j W�f  �M����ܭ �D��E�P�I�I�ѡD�j j��@�@�M�h��Q�СD��M�Q�@�@�Ѓ���j ��� ��_^[��]� _^3�[��]� �������������U���SV��u��^� �E��V� �Ѕ�t7�D�h-� R�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3��u�E��P�e  j �vP���  �oE�����u�� �D�j�vP�@����@V�СD��M�VQ�@�@�Ѓ����u�ŭ �M���j �	� �D��E�P�I�I�у���^[��]� ����������U���<SV��W�]��m� ���}��t:�D�h-� W�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E����3��u�j�Eċ�P�T  �sP���~e  �]����te��I �D����   �΋@��=�� u3�D�V�@@�@,�ЋD����ЋA��j Wh�  �@l��;���   �E����pP��T ����u��u��M�j �vP�   �D��ˋ��   �@��=G  tu=�� uc�D��ˋ��   �@x���oEă����D����u�@j�vP��@����V�СD�VW�@�@�ЋM���hմ �$� ���}�l3�_^[��]� �D��ˋ��   �@x���oEă����D����u�@j�vP��@����V�СD�VW�@�@�ЋM���h�� 趫 ���E��t��E�ύ4��E��P�zV fn΃���ɋ���@�X��X���f���-[ �D�W�@@�@,�ЋD������}�Q��Sh�  �Rp�ҋD��M�j hS  �B�IT���   �ЋM���E��P��U fn΋����� �\��E��@�D��\�����   �E��E܋@��=G  ��   =�� ��  ��  ���$    �j �E��E�    PV�M��E�    �! P����� �M��# �D��M�Q���   �@8�Ѓ���t7�u��oEԃ���SV�u� ������E�� �Xh��E��E���D���j V�@�@0�СD��M�Q���   � ��F�����  �L����E_^[��]� 3����$    ��I V�E�    �E�    ��������M���E�j PW�  P��� � �M��" �D��M�Q���   �@8�Ѓ���td�ƃ�tp��tk��tf�D��MjW�@�@0���u��oEԃ���V� �"�����PS�u�����E�� �Xh��E��E���D��Mj W�@�@0�СD��M�Q���   � ��F���������E_^[��]� ��������������������������VW��跭 ����t5�D�h-� V�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3�V�wP����  j ���������_^�   �������������U���SVW���@� ���}��t5�D�h-� W�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��sP�ȉE���`  ����t9j ���Q ���sP��t�P �M���j�u�V�   ����}P ����uʋ}��D����   ���   ��WP�E��Gw���u�M����	 Pj Vh+� �F ���M��  �D��M�Q���   ���   �Ѓ���j �� _^[��]�������U���S�]V�uWVS�	  �D��]S�@@�@,�ЋD������Q��jh�  �R0�ҋD����   �M�@��-�� tx��t	��&��   ��tKj Sj(���� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ѓ��D���j h�  �@�@p���   �D���j Vh�  �@�@l�ЋȉM��tn��tNj Qj-���Z� �D��M�Q�@�@�СD��M�j j�hض�@Q�@�СD��M�Q�@�@�ЋM���D����   �@L�ЍEP�Q ����tKj Sj-���� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ѓ��D��M���   �@L�ЍEP��� ���} tj j hlcrd�:� ��_^[��]� ��������������U���SVW�}�ى]�����  �E��tF����� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ�W�ˉ}��]  �؅�tW���M �M���j �uS�q����ޅ�u�]��K��t7�D����   �@X�Ћ���t!;�u��� w ����u��jV���ހ ��ujj ���π �]��tKj Wj-���l� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��D��M���   �@L�ЍEP�A� ����tF���� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ�j j hlcrd�v� ��_^[��]� ����������U��E0�����wQ�$��3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø
   ]Ã��]Ë�7;BIPW�^ls��zeU��E������I�  �$��3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø
   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø    ]ø!   ]ø"   ]ø#   ]ø$   ]ø%   ]ø&   ]ø'   ]ø(   ]ø)   ]ø*   ]ø+   ]ø,   ]ø-   ]ø.   ]ø/   ]ø0   ]ø1   ]ø2   ]ø3   ]ø4   ]ø5   ]ø6   ]ø7   ]ø8   ]ø9   ]ø:   ]ø;   ]ø<   ]ø=   ]ø>   ]ø?   ]ø@   ]øA   ]øB   ]øC   ]øD   ]øE   ]øF   ]øG   ]øH   ]Ã��]�Rn����,3�:AHOry�����������!(/|�V]�����6=��u�dk����DK����Y`g����	�%������������U��E������Iww����$����  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]Ã��]�{C�Q<X_f5mt�.�J�  				



		

 		

   ����������U��W�}��tM�D��IV���   �@X�Ћ���t2S�]��$    ���iH ;�ujSj ���L j ���PF ����u�[^_]� ���U���SVW�}�M����*H ���B  j ���G ���1  j ���(G �E����  �]3�V���G ��t[��tKj Wj*���̜ �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ�jj V���QK F��c|��M��Ej PW�E    �E�����^� ������   �d$ ��tKj Vj*���@� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ѓ�j�u����u��J �E�M�@P�E�EPW�E�����֠ ����u�_^[��]� �������U���,SV�u�M�W����  �D��I���   �@X�Ћ�����  �]���F ;��a  j ���F ���P  ���rF ���A  j ����E ���0  j ���pE �E���  3��I V���XE ��t[��tKj Wj*���� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ�jj V���I F��c|��M��Ej PW�E�    �E����覟 ������   ��tKj Vj*��茚 �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ѓ�j�u���u�I �E��M�@P�E��EPW�E�����"� ����u��uj ��� C �����}���_^[��]� �������������U���pVW���P �  �D��GH�OTh�   �@hP  �E؋��   �ЋOTj hQ  fn��D�����@���   �E��ЋOTjhN  fn��D�����@���   �E��ЋD����OTjhO  �R���   ���o_(��3��oG8��W�f(�f(��\O0�\�D��E��M��E�\��E��E�]��\��E��E��U��M���E�f.���]�\��   ��U�\��   ��DzW�fE��U��]���^��^��]��U��U��]��oE���   ����  ���   �X����   ���   �X����   ݇�   �E��ku �]�݇�   �E��Zu fnU��]��o��   ���f(�fTP�f/��]��E��U�w�E��\�f/�w�E��F�E����X�W��^E�f/��E��E��$v�ۑ �贐 �U����]��E��YE��]�f(��E�fTP�f/�w�E��\�f/�w�E��A�E����X�W��^E�f/��E��E��$v�c� ��<� �]��E؃��YE苏�   �E�P�E���B �U�W��M��\�\H�X���X���U��E��E��E��M��E��E��]��E��E��E��U��U��]�f.ܟ��Dzf.ԟ��D��   �o� �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��wP���O  ��3��E���tej ����@ ��t;�E���P��A �M����E����XM��XE؋�f��M���F �E��wP����> ����u��}�u������_^��]� U���  ��3ŉE��EV��E�W�~ �2  脛 �ȅ�t6�D�h-� Q�@L���   �Ћȃ���t�D�j Q�@@�@8�Ѓ����3��E���u���H;  �E�����  ����i �M�������P�]��Ti �u����zN  (p���p����D���f�p���Q����������E��BhW  Q�N���   �}��Ѝ�p���QhX  �o ������Q�N�������~@�D�fօ����( �f�p���W��E��@���   ���U����o �������~@fօ����(��YP�f/���E��E��$v�f� ��?� �N���]��E��\�jhY  �,��E��D��@���   �ЋN�EčE�P�E�P�E�Ph�  �� fnE��E��������NP�E�P�E�P�^�h�  ������fnE�����^�������fnE�����^��������/� fnE��������^���p���fnE�����^���x���fnE�����^��E�����  �I �D�j W�@@�@8�Ѓ��E�3����W�R\�҅��z  �M�W�== �E����f  �������W�u�P��v  �jc�u�� �\�������`����@��t����\�������`���P�M���h�����h����E��v  ��l����]��� �\������U��=���e��\��� ����@�2   �\������������ ����W���(���������������������d����\��f(���H����\��]��U�fTP��Y���,ȃ�2Lȋ���fn������ ����� �����0�����$�����4�����(�����8�����,�����<���fn������@�����@����������D����������H����������L���������}�un��0����X��Y��E���8����X��Y��E�������X��Y��E�������X��Y��E�f(��Y��E�f(��Y��E�}�\�E��\�M�f(�f(��\��\��Y5���Y-���X��X��Y��Y���P�����X�����   9E��   9M��   9}u|�N������P�� �E��E��M����YE�j�u��YM�P���D$�$�%  �o�p���j ���ă�� �E�f�@���o������ �~������  �U ��t	����   9E$��   9M,u}9}(ux�N������P��� �E��M��E��YM��YE��� t*H�o����NPPj�E�P���D$�$�K� �L����,E�NP�,E�P�,�P�,�P�X� �)���j ���9 �N����   h�  �� �E��M��E��YM��YE��� t#Hu>�NPPj�E�P���D$�$��� ��,E�NP�,E�P�,�P�,�P��� �N������P������P������Ph�  �6� �o�p���j ���ă�� �E�f�@���o������ �������   ������P�� �E��M��E��YM��YE��� t#Hu>�NPPj�E�P���D$�$�� ��,E�NP�,E�P�,�P�,�P�� �o�p���j ���ă�� �E�f�@���o������ �~������u�f�@���o�P�������� �\  �E�G��c�g����u��M��6 ���}ȅ��7����M�_3�^�{j ��]�, �����U���@W���O����  V�v� �O�E��� �M�E���a �D��Oh�   hP  �B�]苀�   �ЋOj hQ  fn��D�����@�YE苀�   �E��ЋMfn��E����P�YE��E���` �Oh�  ��H�YU��YM�fW`��U�fW`��M��� �u��u��OVj j ��� �O�E�W�PfE��E��� �,E�O�u�Pj P�k� �,E��OPVPj �Y� �Oh�  �� �E��M��\��E�f/��r4�u��O�,�VPj P�� �E��M��\�f/���E�sҋu��E��X�fn�����E�f/�r0�u��O�,�Pj P��� �E��XE�fn�����E�f/�s��E��M��\�f/���E�r0���O�,�PVPj �� �E��M��\�f/���E�s��E��X�fnM�����E�f/�r6��I �O�,�PVPj �/� �E��E��XE�fn�����E�f/�sϋOj�u� �O�E�W�h�  PfE��E��7� �D��M�Q�@�@�СD��M�j j�hl��@Q�@���E����X��Oj �,��E��X0�P�,�P�E�P�'� �D��M�Q�@�@�Ѓ�^_��]� �����������U��V��~ ��   W��� 3�9~u9~t�   h  �h�  ���� �u���u�u�u�C� �D��5���@�@�Ѓ�����   �N0�F,h   QP�v(�v$QPj j �5�����/� ��tdh�  ���� �F,��j HPj j �� �F0��HPj j j �� h�  ����� �N0�F,IQHPQj ���{� �F0�N,HIPQj Q���g� _^]� �U���XSV��W�E���� �]�ËM+��u�}P��+�PQ�M�W�}� �M�j�� �M�h�  �v� S�]���V�uW�6� �{P tv軎 �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��H�sP��t#�D����   �@X�Ѕ�t;�t����[ ��u��CP    �CP����   j���� ���+���P�y� ( ��+���P���ă�� �X�f�@��(p������ V���f�@�D��@�@�СD�j j�h���@V�@�Ѓ��K�  _^[��]� P�K �2����A���sP�K�C�O����o��   ���   ���̃���A���o��   ���   �sP��A�K�����sP�K�  �sP�K�J  �oCp���K�ă�� ���s\�oC`�sP� ��  �o�  �o�   �E��o�   f~��E��~�0  �E��M���tR�}� �Kth�  �a� �(���E�fE�PW��E��"� �,E��KP�,E�P�,E�P�,E�P��� _^[��]� ���������S�܃������U�k�l$���  VW���}� ��  �>� �ȅ�t;�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ���4����
ǅ4���    �K�Z �s���@���Pݝh����h  ��@����������Y���KP�E���H����Y���E��1 �K� �\E��E��@�������\E�P��p����Y �D��Oj hT  �@���   �Ѓ��E	   fn�����Y�h���f/���E��E��$v�^ ��7~ ��h������Y0����]�f/���E��E��$v�$ ���} �E���Y�����]�f/���E��E��$�E�v��~ ���} ��h������YP���ݝP���f/���E��E��$v�~ ��} �s����ݝ`����0 (����x����D�f�x���Q����������E��E��Bh^  Q�O���   ��j V�o �������������~@�D��E؋@@�@8��������O����fW`�U�j�]��E��U��M���X]���X�p����u��]��U��7� ��h����� ����E�f��Y��� ����E��Y�������@���fY������Y �K�$. �� �������������������� �����t[�O����   h�  �� ������X�����o� ����O�,�f(��X����P�,�P�,����P�,�P�� �P���ϋă� �}� t( �� �H��W�� f�@��(�f�� ��f��@��  �o� �������������������X���X���\=��\-�(0��O�]���p����m���x����h�f�E��� �����ta��x���P�T� �E��XE��o� ����O�,�f(��X�p���P�,�P�,E�P�,�P�	� �o� ����]��m���p����}� f(��E�f(�O�X��Y���X���W��X��u�(��\�(��X��u���8���t( ���x����X�f�M��( ��H���x���f�E���ta��x���P�d� �E��X�8����O�,���X����XE�P�,�P�,E�P�,�X���P�� ��p����m��]��o� ����,U��,�R����f��E��E��X��f���@����,�(�f��,ȉ�<�����<����,�Q�M��O)E�P��\����� �������Q���PP�}� �������O�r  �h��������\��������\��\��Y��Y��Y��X��X��X�������f֝����f���������������tN������P�� �E��XE�O�,���@����XE�P�,�P�u���\������ �������o������,�`���j ���ă���@����XM�( ��e��Xe���\�P���f�X��Q���e���� �X�f�@��f����  �K�E�P��, �D��ЋA�ʋ@<�ЋD�����E�P�I�I�у�����   �-�������������������\��h��\��e؃�( ��\�����X��Y��Y��Y���@����X��X�P����X�f�H���X�f���`����X���f�`�,��E�P��fЋ���?  ����U��,E�j(0��Y�P(`��X�@����,�P���ă�� �h�f�@���f�X��  f֝�����o�������������tN������P��� �E��XE�O�,���@����XE�P�,�P�u���\����� �������o������,�`���j ���ă���@����XM�(`��e��Xe���\�P���f�X��Q���e���� ���f�@��f���  �K�E�P��* �D��ЋA�ʋ@<�ЋD�����E�P�I�I�у�����   �o���������������e�(�f(�f��Y�f(ă��Y��Y���@����X�P���f��f�@����`����X���(f�`�,��E�P��fЋ���=	  �U�W��Y��j�,E��X�@���( �P�,�P���ă�� f�@������f�@�K�U��0& �D�������IV�I�ыD�VW�A�@�Ћ}�����  fnE��O���j�XE��,��u���� �K�&) ����  �D��Ojh_  �@���   ��@������+��fn�����Y�h����E��E��$�'u �,E����O��p����X��Pݝh����,�P�,� ����u�P�?� �,�h������oE�fn�����\��M��,�fn�����Y���E��E��$�t �]��,E؋Kj Qfn�����X�@����,�fn�����E��D��@@�E��XE��@8�,��Ѓ���t;�H0��t4�}� �  �   EU�P�,�h���jZjZj j PPVRQ�O�� �?�O������W�Pf������������>� �,�h����U��P�
�OPVR�� �E��Y��XE��XE��,��u��D��Oj h]  �@���   �Ѕ���   �K�E�P�& �D��M��@�@<�Ѕ���   �,E�Ofn����P��<����,��E�P��\����� �E��XE�j�,�P�,E�P���ă��}� ��Vt(`�����(������f�@�D��@�@�СD��M�VQ�@�@�Ѓ����  �E��XE��,��u��D��M�Q�@�@�Ѓ��K������P��$ �D��������@�@<�Ѕ���   �,E�Ofn����P��<����,��E�P��\����� �E��XE�j�,�P�,E�P���ă��}� ��Vt(`�����(������f�@�D��@�@�СD�������VQ�@�@�Ѓ����  �E��XE��,��u�u��u����E�    ��@d�Ѕ���  3ɋQ�΋@\�Ѕ���  �,E�OfnE����P��<����,��E�P��\����� �}� ��u��,  �M�Q���PX(P��O���������fօ������tHh�  ������P�p� �E��XEȋOj�,���@����XE�P�X0��,�P�E�P�� �D��M�Q�@�@����@������X�P����K�u��������E��XE��E��  (0����o��������@P���ă�� �h�f�@��( �� �X�f�@�,�`����E�P��fȋ����  �9  �M�Q���PX(`��O���������fօ������tHh�  ������P�D� �E��XEȋOj�,���@����XE�P�X0��,�P�E�P�]� �D��M�Q�@�@����@���������X�P�������u��@`������Q�E����XE��E����u��K���r (0����o��������@P���ă�� �h�f�@���o� �~Ff�@�,�`����E�P��fȋ���  �u��E��XE��,��E����E��@d�ЋM�;��%�����΋@T�Ѕ���  �,E�O��p����X��fnM�P����,�P�,�P�,� ���P��� ��4����E�j P�s�Ty �ȋE������fn��}� �M����t~(0�3�( ����o� ������U��X�p���P���Xԋă��\�P���� �h�f�@���X�f��f�@�,�`���P������   �o� ���������jc�X�p���Q�@`���\�P����� ����E��X��E���(0�3�9M����o� �����Q���̃�����h�f�A�o� �~Bf�@�,�`����E�P��fȋ������  �O�Y� �OP�0� �OPj j �c� �D�������Q�@�@�Ѓ�_^��]��[� �U���8fnEW����V�����Y��f/��E��E��$v�l ��k �M�   �U���]��,E�W�;�L��Nfn�����\��\��oE4�X��X��E��~ED�M��U�f�E؅�tL�E�P苼 fnM��ɋNf(��XE��,�f(��XE�P�,�P�,E�P�,E�P�B� �M��U��X���X���oE�N�M�fnM�U�����E��~E,(�f�E��\��\��U��M��t;�E�P�� �E��XE��N�,��E��XE�P�,�P�,E�P�,E�P袿 ^��]�D �����������U������tfnE���SVW���L$H�Y��f/���D$P�D$P�$v� k ���i �m�   �\$P�,L$P��f(�;�LȉL$Dfn�����\��,�f(��Xŉ|$0fn����f/��7  � ��}�����]׉T$4f(��\��,�f(��XÉ\$(fn����f/���  �4I�]����ˉL$,�I W��Yڋ��D$<   �D$Hf(��YD$8�\$P�D$`�fnȋ���ɻ   �\��Y��L$X�I fn�����\��Y��X���g fn����f/�w.�}L tf(��\ �f/�w�T$H�X���T$H��T$H�L$XG�\$PKu��D$8�D$`@�L$<�L$,�D$8�X����^P�f.�����D{v�M�D$h�\M4�L$@P�YʋI�XM4�L$l�M$�\M<�Y��XM<�L$t�M,�\MD�Y��XMD�L$|�f� �|$0�\$(�D$@WSW�HS�>� ��\$(�|$0�D$DC�]�L$,� ����m�T$4fn����\$(�L$,fn����f(��X�f/��H�����Gf(��Xŉ|$0���T$4fn����f/������_^[��]�H �������U���4S�ى]��{ �*  �%t �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3�VW�}��W�K'  ������   ���E�VP���P  �E܍E��Y����P�E��E��Y���E�� �C(�U��M�� �X�\e��\]��k�Y��Y��Y��Y��C�X�f/�w6�X�f/�w,�S�C �X�f/�w�]��X�f/�wWV��������]�W���< �����2���_^[��]� ���������U���  ��3ŉE�V�uW��� �<  ��u��r P�0��������  �����  ���RA ��������Pݝ������@ �Oj�4� �������������$hp�P�I ��W�j jjh�  ���ă���� Vf�@�D��@�@�СD�������j j�Q�@V�@�Ѓ����   ���������������$h|�P�H �O��j �� ��W�Pjh�  ���ă���� Vf�@�D��@�@�СD�������j j�Q�@V�@�Ѓ����  �M�_3�^�H ��]� ��������������U��V��N��t;�E(P�ڵ �E �XE�N�,��E�XEP�,�P�,EP�,EP蘹 ^]�8 ���U��Q�} W����   �M �Ef/�vf(��f(��](�,��Uf/ډE�vf(��f(�f/��,ĉEw(�f/�SV�,�w(ӋOh�  �,��D� �E�OPSP�u��Ӹ �OVS�uS�Ÿ �OV�u�VS跸 �u�E��OPVP覸 ^[_��]�( �������������U��E�U�� t,HuI�E�IPPjR���D$�E�$�*� ]� �,B(�IP�,B P�,EP�,EP�6� ]� ��U��V��N��t#h�  �EP�e� �u8�N�E�u4�u0P蠸 �D��MQ�@�@�Ѓ�^]�4 �������U��S�ًK��teVWh�  �E0P�� �������uP�EL�K�P�EH�P�EP�B� F��~�G��~֋K�Eh�  P�մ �uP�K�E�uL�uHP�� _^�D��MQ�@�@�Ѓ�[]�L �����U��S�ًK��teVWh�  �u0�d� ��������u<�E8�K�P�E4�P�EP買 F��~�G��~֋K�Eh�  P�E� �u<�K�E�u8�u4P耷 _^�D��MQ�@�@�Ѓ�[]�8 �����U���SVW���pn ��ˉE��Rl������   �u�E�j P�u�E�   �u��1�  ���M�P�E� P��證 �M��E� �D��M�Q���   � �Ѓ���tm��!���D���j hS  �A�ʋ��   �ЋK���E��P�� �u�fn��������\��@�\�����uW�sf���!����� jj���� j �y ��_^[��]� U���SVW���pm ��ˉE��Rl������   �u�E�j P�u�M��E�   �u��N� P��趈 �M��N� �D��M�Q���   � �Ѓ���tm�� ���D���j hS  �A�ʋ��   �ЋK���E��P�� �u�fn��������\��@�\����W�u�sf���J����� jj���� j �x ��_^[��]� ���������j j h�� �Rx ���   � �������j j hɴ �2x ���   � �������j j h�� �x ���   � �������j j h�� ��w ���   � �������j j h�� ��w ���   � �������j j h�� �w ���   � �������j j hô �w ���   � �������j j h�� �rw ���   � �������j j h�� �Rw ���   � �������j j h�� �2w ���   � �������h'� � ���   � �����������j j hǴ ��v ���   � �������j j h�� ��v ���   � �������j j h´ �v ���   � �������j j hƴ �v ���   � �������j j hĴ �rv ���   � �������j j hŴ �Rv ���   � �������j j hl� �2v ���   � �������j j ho� �v ���   � �������j j hf� ��u ���   � �������j j hy� ��u ���   � �������j j hg� �u ���   � �������j j h�� �u ���   � �������j j hm� �ru ���   � �������j j hh� �Ru ���   � �������j j h�� �2u ���   � �������j j hp� �u ���   � �������j j h�� ��t ���   � �������j j hq� ��t ���   � �������j j hr� �t ���   � �������j j hs� �t ���   � �������j j hi� �rt ���   � �������j j h�� �Rt ���   � �������j j hj� �2t ���   � �������j j h{� �t ���   � �������j j hz� ��s ���   � �������j j h�� ��s ���   � �������j j h}� �s ���   � �������j j hx� �s ���   � �������j j hk� �rs ���   � �������j j ht� �Rs ���   � �������j j h�� �2s ���   � �������j j hu� �s ���   � �������j j hw� ��r ���   � �������j j h�� ��r ���   � �������j j h�� �r ���   � �������j j h�� �r ���   � �������j j hn� �rr ���   � �������j j hd� �Rr ���   � �������j j h~� �2r ���   � �������j j h|� �r ���   � �������j j he� ��q ���   � �������j j h�� ��q ���   � �������j j hv� �q ���   � �������j j h� �q ���   � �������j h,  h�  j�j�h&� j���Ѷ � ��������������U���PVW���M��t4�D�h-� Q�@L���   �Ћȃ���t�D�j Q�@@�@8�Ѓ��3��H����  �D����   �@X�Ћ�����  �d$ ���2 ��u���n2 ����u�_�F^��]� ���b  ���X  j���������"  �w���4 ���  �D��M�SQ�@�@�СD��M�j j�hp��@Q�@�СD��M�Q�@�@�СD��M�j j�ht��@Q�@�Ѓ�(�E�j$P�G@P�E�P�Y{  P�E�P�E�P�{W����P�E�P�nW����P�k ���MСD�Q�Ë@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���[�;  �w����5 _�   ^��]� �w���]3 ���w��t#�?6 j j h,� �Qo ���   _^��]� �7 �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E�j@P�G@P�E�P�z  P�E�P�E�P�1V����P�E�P�$V����P�Kj �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��@�@�M�Q�Ѓ�_�   ^��]� ������Vj h,  h�  j�j�h�� j��萳 ����tj j h�� �n ����^� ���U���HSVW���b �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3�(@����sPfE�3�(p�fE��  �]Ћ�����   �E��E��E��E��E��]��E�j ���$ ��tN�E���P�U �M��E�f/�v�M��E��U�f/�v�E�f/M�v�M�f/E�v�E�G�sP���H ����u��M��U��]��e���e��M��U��\��\��Y���Y���X��X��U��E��E��E��M��E��E��E��E��E��~b���� �M؋˙+���fn�����\��M��ޣ �M����KP�+���fn�������\��oE�f�� �1 j ��蕢 _^[��]���������������� �������������U��} t�M��t�j�]� �����̋IV��t0�D����   �@X�Ћ���t�����y- ��u���>- ����u�3�^Ë�^áD�Q���   �@8�Ѓ������������U��U�A��A�B�B*� �B   �A�B�A �B�   �B)� �B   ]� ��������������U��D���@�@V�uV�@�СD�j j�h���@V�@�ЋE�����g  �$�L�D��M�Q�@�@�СD��M�j j�hȿ�@Q�@�СD��M�VQ�@�@�СD��M�Q�@�@�Ѓ� ��^��]� �D��M�Q�@�@�СD��M�j j�hп�@Q�@�СD��M�VQ�@�@�СD��M�Q�@�@�Ѓ� ��^��]� �D��M�Q�@�@�СD��M�j j�hԿ�@Q�@�СD��M�VQ�@�@�СD��M�Q�@�@�Ѓ� ��^��]� �D��M�Q�@�@�СD��M�j j�hؿ�@Q�@�СD��M�VQ�@�@�ЋD��E�P�I�I�у� ��^��]� ���J�JYK�K�D����   ���   ���������������U���dV��M��FH�E�W�fE���u �E��E�    Pjhsuom���E�    �� ���  �D��M�j hxvpi�@���   �ЉE��M��D�j hyvpi�@���   �ЉE��΍E�P�E�P�\� �} ufnE��u����fnE������   �oF8�of(�E�fnE�(����f��X��E�fnE��U��M�����f/��X��E��E��E��E��E�vf(��E��X�f/�vf(��E�f/�vf(��M��X�f/�v(��
�E��U��]�Wɋuf.ٟ��Dz�M���t ��^��]� �^��^���M��F��t ��^��]� ��������U����D�S�]�M��ˋ��   W�@�Ћ}��P�U� ��u_[��]� �D�VS�@@�@,�ЋD��������   ���   �щE���u3��   �D�S���   �ȋ��   �СD���j h�  �@���   �ЉE�M��E��E�_  P�E�    �E�    �� �u��E���P��� �M������ ��t�D��A3�9M���@0Qj���СD���jh�  �@���   �ЉE�M��E��E�Z  P�E�    �E�    �� �u��E���P�]� �M����� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�V  P�E�    �E�    �� �u��E���P��� �M����� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�S  P�E�    �E�    �#� �u��E���P�u� �M����� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�a  P�E�    �E�    �� �u��E���P�� �M����'� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�U  P�E�    �E�    �;� �u��E���P�� �M����� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�W  P�E�    �E�    ��� �u��E���P�� �M����?� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�X  P�E�    �E�    �S� �u��E���P�� �M������ ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�Y  P�E�    �E�    ��� �u��E���P�1� �M����W� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�\  P�E�    �E�    �k� �u��E���P�� �M������ ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�]  P�E�    �E�    ��� �u��E���P�I� �M����o� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�R  P�E�    �E�    �� �u��E���P��� �M������ ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�^  P�E�    �E�    �� �u��E���P�a� �M����� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �ЉE�M��E��E�T  P�E�    �E�    �� �u��E���P��� �M����� ��t�D��A3�9M���@0Qj���СD���j h�  �@���   �Ћ��E�`  �E��E�    P�M��E�    �(� �u��E���P�z� �M����� ��t�D��A3Ʌ����@0Qj���Ћuj ��U` �M���VW�u�ew ���D��E�P���   ���   �у���^_[��]� �������������U��Q�D�V�u�M��@@�@,�ЋM����j ��� ����  tuItM��t�u�M��u�u�u�u�  ^��]� �D���j h�  �@���   ��3Ƀ�^������]� �D���j h�  �@���   ����^�@��]� �D���j h�  �@���   �Ѕ�t&�D���j h�  �@���   �Ѕ�t	3�^��]� �   ^��]� �����������U��Q�D�V�u�M��@@�@,�ЋM����j ��� ����  t,��t�u�M��u�u�u�u� ^��]� j h�  �j h�  �D��΋@���   ��^��]� ���U��Q�D�V�u�M��@@�@,�ЋM����j �i� ����  t:��t,��t�u�M��u�u�u�u�~ ^��]� j h�  �j h�  �j h�  �D��΋@���   ��^��]� �����U��Q�D�S�u�M��@@�@,�ЋM����j ��� �8�  t�u�M��u�u�u�u�� [��]� �D���j h�  �@���   ��3Ƀ�[������]� ���������U��Q�D�V�u�M��@@�@,�ЋM����j �Y� ����  t!It�u�M��u�u�u�u�u ^��]� �D���j h�  �@���   ��^��]� ��������������U��Q�D�S�u�M��@@�@,�ЋM����j ��� �8�  t�u�M��u�u�u�u�� [��]� �D���j h�  �@���   ��3Ƀ�[������]� ���������U��Q�D�V�u�M��@@�@,�ЋM����j �Y� ����������   �$�tZ�D���j h�  �@���   �Ѓ�tc�D���j h�  �@���   �Ѓ�tE�D���j h�  �@���   �Ѓ�t'�D���j h�  �@���   �Ѓ�t	3�^��]� �   ^��]� �D���j h�  �@���   ��3Ƀ�^������]� �D���j h�  �@���   �Ѕ�t��D���j h�  �@���   �Ѓ��'����u�M��u�u�u�u�u ^��]� ��_Y�Y�YZ������������U��Q�D�S�u�M��@@�@,�ЋM����j ��� �8�  t�u�M��u�u�u�u�
 [��]� �D���j h�  �@���   ��[��]� ���U��Q�D�V�u�M��@@�@,�ЋM����j �y� ����  |`���  ~2���  uP�D���j h�  �@���   ��3Ƀ�^������]� �D���j h�  �@���   ����^��؋�]� �u�M��u�u�u�u�8 ^��]� �U���V�q8�E��  V�E��E�    P�ު ��u�V�E�   �    �B    �    �D��E�j ���   �E�PR�I�ыD��E�P���   �	�у���^��]� ��������������U���V�u葨 �D����E�P�I�I�ыD��A�M�QV�@�СD��M����@�@<�Ћu���D�V�@�@t2�СD�V�H�E�P�I�ыD��E�P�I�I�у���^��]� �СD�j j�hL��HV�I�ыD��E�P�I�I�у���^��]� �����������U��D��IW�}���   �@X��u��_]� V�Ћ���t�d$ ���� ;�tj ���|� ����u�^3�_]� ��^_]� �����̋I��u3�áD����   �@X�������̸�� �����������U��D��IW�}���   �@\��u��_]� V�Ћ���t�d$ ����� ;�tj ���|� ����u�^3�_]� ��^_]� �����̡D�Q���   �@8�Ѓ�������������VW���wK �D����v�I@�I,�у���Wh�  ��d _^��U��E�Q,��E�I0��   ]� ����U���@V����(��M����E�fE�P�P��E���2���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V�t���(���M����E�fE�P����E��M2���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V�����(���M����E�fE�P����E��1���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V�4���(@��M����E�fE�P����E��1���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V����(���M����E�fE�P�H��E��m0���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ����U���@V�����(���M����E�fE�P�p��E���/���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ����U��E(�� �x��@]� ��������������̸   ����������̸   ����������̸   ����������̸   ����������̸
   ����������̸   ����������̸I   �����������U���u�u�� �E]� �����������U��U�B���	w�E( � �@]� R�u� �E]� ������������U��E��u%�E��������@�H]� P�u�7 �E]� U��E��u�E( � �@]� P�u� �E]� U��E( � �@]� �������U��E��
}�E( � �@]� P�u� �E]� ���������������U��E��}�E( � �@]� P�u�v �E]� ���������������U��SVW��3��   ��KV�� ��E�F��
~�M��t�G;�~��ct	_^3�[]� _^�   []� ����U��E��x��~��cu	�   ]� 3�]� �������������U��E�� tAHt��bt93�]� �D��q�@@�@,�ЋD����ЋA��j h8  ���   ��]� �   ]� �����������U��3��}c��]� U��D��q�@@�@,�ЋЃ��E��
�G  �$��f�D�j h�  �A�ʋ��   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� �D���j h�  �@���   ��]� 3�]� �I [eye�e�e�e�e
f'fDfaf~fU��E��cwJ��8g�$�,g�D��q�@@�@,�ЋD����ЋA��j h8  ���   ��]� �   ]� 3�]� �g�f%g   ����U��3�9E��]� �U��E��t��ct3�]� �   ]� ��U��SVW�����3��I �KV�� ��E�F��
|�M�G_^[;�~��ct3�]� �   ]� �����������U��E��x��~��cu	�   ]� 3�]� �������������U��D�V�q�@@�@,�Ћ����E��H�~  �$��t�D�j h/  �A�΋��   �Ѕ��U  j h�  �)  �D���j h0  �@���   �Ѕ��(  j h�  ��  �D���j h  �@���   �Ѕ���  j h�  ��  �D���j h  �@���   �Ѕ���  j h�  �  �D���j h  �@���   �Ѕ���  j h�  �u  �D���j hG  �@���   �Ѕ��t  j h�  �H  �D���j hH  �@���   �Ѕ��G  j h�  �  �D���j hI  �@���   �Ѕ��  j h�  ��
  �D���j h  �@���   �Ѕ���
  j h�  ��
  �D���j hK  �@���   �Ѕ���
  j h�  �
  �D���j hL  �@���   �Ѕ���
  j h�  �g
  �D���j hM  �@���   �Ѕ��f
  j h�  �:
  �D���j h  �@���   �Ѕ��9
  j h�  �
  �D���j h  �@���   �Ѕ��
  j h�  ��	  �D���j h  �@���   �Ѕ���	  j h�  �	  �D���j h  �@���   �Ѕ���	  j h�  �	  �D���j h  �@���   �Ѕ���	  j h�  �Y	  �D���j h  �@���   �Ѕ��X	  j h�  �,	  �D���j h%  �@���   �Ѕ��+	  j h�  ��  �D���j h&  �@���   �Ѕ���  j h�  ��  �D���j h3  �@���   �Ѕ���  j h�  �  �D���j h4  �@���   �Ѕ���  j h�  �x  �D���j h  �@���   �Ѕ��w  j h�  �K  �D���j h  �@���   �Ѕ��J  j h�  �  �D���j h  �@���   �Ѕ��  j h�  ��  �D���j h  �@���   �Ѕ���  j h�  ��  �D���j h'  �@���   �Ѕ���  j h�  �  �D���j h(  �@���   �Ѕ���  j h�  �j  �D���j h5  �@���   �Ѕ��i  j h�  �=  �D���j h6  �@���   �Ѕ��<  j h�  �  �D���j h  �@���   �Ѕ��  j h�  ��  �D���j h  �@���   �Ѕ���  j h�  �  �D���j h  �@���   �Ѕ���  j h�  �  �D���j h  �@���   �Ѕ���  j h�  �\  �D���j h)  �@���   �Ѕ��[  j h�  �/  �D���j h*  �@���   �Ѕ��.  j h�  �  �D���j h7  �@���   �Ѕ��  j h�  ��  �D���j h8  �@���   �Ѕ���  j h�  �  �D���j h  �@���   �Ѕ���  j h�  �{  �D���j h  �@���   �Ѕ��z  j h�  �N  �D���j h  �@���   �Ѕ��M  j h�  �!  �D���j h  �@���   �Ѕ��   j h�  ��  �D���j h+  �@���   �Ѕ���  j h�  ��  �D���j h,  �@���   �Ѕ���  j h�  �  �D���j h9  �@���   �Ѕ���  j h�  �m  �D���j h:  �@���   �Ѕ��l  j h�  �@  �D���j h  �@���   �Ѕ��?  j h�  �  �D���j h   �@���   �Ѕ��  j h�  ��  �D���j h!  �@���   �Ѕ���  j h�  �  �D���j h"  �@���   �Ѕ���  j h�  �  �D���j h-  �@���   �Ѕ���  j h�  �_  �D���j h.  �@���   �Ѕ��^  j h�  �2  �D���j h;  �@���   �Ѕ��1  j h�  �  �D���j h<  �@���   �Ѕ��  j h�  ��  �D���j h  �@���   �Ѕ���  j h�  �  �D���j hA  �@���   �Ѕ���  j h�  �~  �D���j hB  �@���   �Ѕ��}  j h�  �Q  �D���j hC  �@���   �Ѕ��P  j h�  �$  �D���j h  �@���   �Ѕ��#  j h�  ��  �D���j h1  �@���   �Ѕ���  j h�  ��  �D���j h#  �@���   �Ѕ���  j h�  �  �D���j hD  �@���   �Ѕ���  j h�  �p  �D���j hE  �@���   �Ѕ��o  j h�  �C  �D���j hF  �@���   �Ѕ��B  j h�  �  �D���j h$  �@���   �Ѕ��  j h�  ��   �D���j h2  �@���   �Ѕ���   j h�  �   �D���j h  �@���   �Ѕ���   j h�  �   �D���j h
  �@���   �Ѕ���   j h�  �e�D���j hJ  �@���   �Ѕ�thj h�  �?j h=  �j h>  �j h?  �j h@  �D��΋@���   �Ѕ�t'j h�  �D��΋@���   �Ѕ�t
�   ^]� 3�^]� ��|h�h�hi1i^i�i�i�ij?jlj�j�j�j kMkzk�k�kl.l[l�l�l�lm<mim�m�m�mnJnwn�n�n�n+oXo�o�o�op9pfp�p�p�pqGqtq�q�q�q(rUr�r�r�r	s6scs�s�s�stDtnt�t�t�t�tU��� V�u�F���	wu�D��M�Q�@�@�СD��M�j j�h���@Q�@�ЍF�P�E�P�VJ  �uP�E�PV�x&���D��H�E�P�I�ыD��E�P�I�I�у�0��^��]� ��u5�D��uV�@�@�ЋD�j j�h0��IV�I�у���^��]� V�uV�V� ��^��]� �������������U��U��V�u�� t*HtRV�%� ��^]� �D�V�@�@��j j�hl���D�V�@�@��j j�hd��D�V�I�I�у���^]� �����U��EV�u��u0�D�V�@�@�ЋD�j j�h���IV�I�у���^]� PV�� ��^]� ����U��EV�u��tPV�k� ��^]� �D�V�@�@�ЋD�j j�h���IV�I�у���^]� ����U��U��V�u�� tFHt*HtRV�� ��^]� �D�V�@�@��j j�h,��0�D�V�@�@��j j�h`���D�V�@�@��j j�hX��D�V�I�I�у���^]� ���������U��U��V�u�� t*HtRV�� ��^]� �D�V�@�@��j j�h,���D�V�@�@��j j�h���D�V�I�I�у���^]� �����U��U��V�u�� tFHt*HtRV�� ��^]� �D�V�@�@��j j�h,��0�D�V�@�@��j j�hl���D�V�@�@��j j�hd��D�V�I�I�у���^]� ���������U��EV��
�  �$��z�Mj h���z���E^]� �Mj h���c���E^]� �Mj h���L���E^]� �Mj h̸�5���E^]� �Mj hܸ����E^]� �Mj h�����E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h�����E^]� �Mj h�����E^]� �uPV�� ��^]� �I �y�y�y�yz*zAzXzoz�z�z������������U��EV�u��u0�D�V�@�@�ЋD�j j�h���IV�I�у���^]� PV��� ��^]� ����U��EV�u��tPV��� ��^]� �D�V�@�@�ЋD�j j�h���IV�I�у���^]� ����U���0V�u��
��   �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�VQ�@�@(�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��uV�@�@�СD��M�VQ�@�@�СD���8�΋@�@<�ЋD�j�j��Q�M�QP�΋BL�СD��H�E�P�I�ыD��E�P�I�I�у���^��]� V�uV�� ��^��]� ��������U���u�u�r� �E]� �����������U���0V�u����   �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��H�FP�E�P�A(�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��uV�@�@�СD��M�VQ�@�@�СD���8�΋@�@<�ЋD�j�j��Q�M�QP�΋BL�СD��H�E�P�I�ыD��E��I�IP�у���^��]� V�uV�N� ��^��]� �����U��EV��H��  �$����Mj h������E^]� �Mj h������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h���y���E^]� �Mj h��b���E^]� �Mj h$��K���E^]� �Mj h4��4���E^]� �Mj hH�����E^]� �Mj h\�����E^]� �Mj hp������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h���|���E^]� �Mj h��e���E^]� �Mj h(��N���E^]� �Mj hH��7���E^]� �Mj hh�� ���E^]� �Mj hx��	���E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h�����E^]� �Mj h(�����E^]� �Mj hH��h���E^]� �Mj hX��Q���E^]� �Mj hp��:���E^]� �Mj h���#���E^]� �Mj h������E^]� �Mj h�������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h(�����E^]� �Mj h8�����E^]� �Mj hP�����E^]� �Mj hp��k���E^]� �Mj h���T���E^]� �Mj h���=���E^]� �Mj h���&���E^]� �Mj h������E^]� �Mj h������E^]� �Mj h������E^]� �Mj h0������E^]� �Mj hP�����E^]� �Mj hp�����E^]� �Mj h������E^]� �Mj h���n���E^]� �Mj h���W���E^]� �Mj h���@���E^]� �Mj h���)���E^]� �Mj h�����E^]� �Mj h������E^]� �Mj h0������E^]� �Mj hH������E^]� �Mj h\�����E^]� �Mj hl�����E^]� �Mj h|�����E^]� �Mj h���q���E^]� �Mj h���Z���E^]� �Mj h���C���E^]� �Mj h���,���E^]� �Mj h������E^]� �Mj h�������E^]� �Mj h������E^]� �Mj h(������E^]� �Mj h4�����E^]� �Mj hH�����E^]� �uPV�� ��^]� �~.~E~\~s~�~�~�~�~�~�~+BYp�������(�?�V�m�������ɀ�����%�<�S�j�������Ɓ݁��"�9�P�g�~�����Âڂ���6�M�d�{�������׃���3�J�a�x�������U���(�D�SV���E�    �@Wj�N���   h_  �u���@����+ȡD��j �M��@�NhS  ���   �ЋD�3ۋNShT  �R�E싒�   ��S�u�E	   �E�D��@@�@8�Ћ�����3���Rd��~���W�P\��tC���G�Pd;�|��u����PT���   E١D��M�j h]  �@�I���   �Ћu��t,�E��E�   P����� �D��ЋA�ʋ@<���E���u�E� �E�t�D��M�Q�@�@�Ѓ��}� �   �   ��E��E�P��� �D��ЋA�ʋ@<�ЋD����E�P�Q�R�҃���tG�M� � ��t�U����3�fnE��M�E���_^���[� fn�����@��]� U���X�D�SV���E�    �@Wj�K���   h_  �]��Ћu@����+ȍE��V�M��P������E��E��Y����P�E��E��Y���E��f� �Kj hT  � �\E��E��@�D��\EЋ@�Eȋ��   ��3��E�    SVfnȡD���ɋ@@�Y��@8�XP�f(��M��Y���E�f(��X���E��Ћ����EW��� ��� ��t�E��fn�����XE��E�D��M�j h]  �@�I���   �Ѕ�t,�E��E�   P����� �D��ЋA�ʋ@<���E��u�]�E�t�D��M�Q�@�@�Ѓ�8]t�E��XE��E�E���P�� �D��ЋA�ʋ@<�ЋD����E�P�I�I�у���t�E��XE��E���3��Pd��~*��I ���V�P\���E�t@�E�;u��D؋F�Pd;�|ۃ}c�E�u>�XE��E_^[�\���\E�� �E��XE��XE��\���@��]� �X���M�C��M��XM�_�XE�^[�fn�������YE��X��XE��A��]� ����������̡D�jQ�@�@H�Ѓ�������������̡D�j Q�@�@H�Ѓ��������������U��E�  ��   ]� ����������̸T�����������̸   @� ��������U��UVW����t4�D�h-� R�@L���   �Ћȃ���t�D�j Q�@@�@8�Ѓ��3��H��t.�D����   �@X�Ћ���t����� ��u���� ����u�3��G���u_3�^]� ��t�P����� ��_�%���?   @^]� ����̸�������������U���VW���� �M���g6 �E�P�u�N�u �D��M�j Wheert�@�@l�ЍM���6 _��^��]� ������������U���`�MSVW�o �]��D�S�@�@�СD��MSQ�@�@�Ѓ��E   ����   ���    �D��΋��   �@x�ЋD����E�P�I�I�ыD��A�M�QW�@�СD��MЃ��@S�@x�Ѕ��D�tG���   �΋@(�Ћ��MСD�Q�@�@�Ѓ���u��D��EP�I�I�у���_^[��]� �@�M�Q�@�СD��M�j j�h���@Q�@�СD��M��uQ�@�@(�ЋD����E�P�I�I�ыD��A�M�QW�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�MQ�@�@�СD��M���8�@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�СD��M�Q�@�@�M�Q�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�SQ�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M��EQ�@�@�Ѓ��������������̡D�Q���   �@@�Ѓ�������������U��D��u�u�@�uQ���   �Ѓ�]� ������������U��D����@SVW�}�񋀠   ��j hacpi�Ѓ~P �؉^Xj uj h�� �P& ���   _^[��]� �D����E    �E�    hxvpi�@���   �ЉE�ϡD�j hyvpi�@���   �ЉE��΍E�P�EP�e fnM��fnE����j �������f���E�P�@O  �D���j haqpi�@���   �Ѓ�Ku�M��u�M��t��t��� ��b� j �% ���   _^[��]� ����������U��D�SVW�@�ًMj hacpi���   �ЋD����Mj haqpi�R���   �ҋȋ�у�������cOt�ǽ����   ��x��$�d�����   ����   ����   QQh�� ��$ ���   _^[]� ��xmtD��dt,��vui��te��ua��u]QQh�� �$ ���   _^[]� ���� _^�   []� ��t+��u'��u#QQh�� �[$ ���   _^[]� ���  t	_^3�[]� j j h�� �-$ ���   _^[]� ������Ӑ�<� ��U��D���0�@S�]V���   ��Wj hacpi���Ѓ~P ���~Xu&���%  h���h������T �G�_^[��]� hTCAb�M��E�    �E�    �]0 �M��50 ���Z �D�Phdiem�Q�MЋB4�СD��M�j havem�@�@4�СD���j hxvpi�@���   �ЉE��ˡD�j hyvpi�@���   �ЉE��΍E�P�E�P�b �D���j haqpi�@���   �Ћ؃�tt��to��tj��d�  �D��Mj havpi�@���   ��fnM���fnE���Q�ˋЃ���Q���S���΋����Rf���J  j ����X �  �M��fnM�fnE�QP�Ë΃���P���S�������Wf���|<  j ���X �E��P�vXhsuom� Z ���^  ���    �D��M�j hxvpi�@���   �ЉE��M�D�j hyvpi�@���   �ЉE��΍E�P�E�P�ga �D��M�j haqpi�@���   �ЋD���j havpi�Q�M䋒�   ��fnM���fnE�����ɋ����f�tg��P�ǃ���PW�����vX���C  j ���W �D��M�jhrdem�@�@4�ЍEЋ�P�8X �E��P�vXhsuom�Y ��������Q��P�ǃ���PW�����vX��,F  j ���SW �FX    �MСD�j hrdem�@�@4�ЍEЋ�P��W j ��  ���M��- �M��- _^�   [��]� ��U���V�uV�� �D�V�@@�@,�ЋD������Q��jh�  �R4�ҋD�������A���$h�  �@,�СD���jh9  �@�@4�СD��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M����@Qh<  �΋@8�СD��M�Q�@�@�Ѓ��   ^��]� �����U��V�uV�3� �D�V�@@�@,�ЋD�����Q�$�Q��h�  �R,�ҡD������΋@�$h�  �@,�СD���jh�  �@�@0�СD���j h�  �@�@4�СD�������΋@�$h�  �@,�СD���jh�  �@�@4�и   ^]� ������������U���V�uV�P� �D�V�@@�@,�ЋD������Q��jh�  �R0�ҡD��M�W�fE�Q�E��΋@h�  �@H�СD���jh�  �@�@0��( ��M�D�fE�Q������E��@h�  �@H�СD�������΋@�$h�  �@,�и   ^��]� ����������U���   V�uV�m� �D�V�@@�@,�ЋD������Q��jh�  �R4�ҋD�j h�  �A�΋@4����� �E��u3���   ����M����W��E��E�W��E�Q( ����U��E�    �U��E�    f�M��M��E�f�U��U��Q� �M�E�P�E� �D��M��u�E�    �E�    ���   h!D Q�@\�СD��M����@Qh�  �΋��   �СD��M�Q���   � �Ѓ��   �EP�9� ����^��]� �������������U���V�uV�� �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD�j h�  �A�΋@4�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@Qh<  �΋@8�СD��M�Q�@�@�Ѓ��   ^��]� ���������U���V�uV�P� �D�V�@@�@,�ЋD������Q��jh�  �R4�ҋD���W��A���$h�  �@,�СD���jh�  �@�@0���;� �E��tmj���;� �E��t]�D�P�E�    �E��E�    ���   h�e P�A\�СD��M����@Qh�  �΋��   �СD��M�Q���   � �Ѓ��EP�� ���   ^��]� ���������������U��V�uV�C� �D�V�@@�@,�ЋD������Q��jh�  �R0�ҋD�jh�  �A�΋@0�СD���jh�  �@�@0�СD���j h�  �@�@4�СD���jh�  �@�@4�СD���jh�  �@�@4�и   ^]� U���V�uV萿 �D�V�@@�@,�Ѓ����Ț �E��tmj���Ȝ �E��t]�D�P�E�    �E��E�    ���   h�e P�A\�СD��M����@Qh�  �΋��   �СD��M�Q���   � �Ѓ��D�������΋@�$h�  �@,�ЍEP�W� ���   ^��]� ��������U��V�uV賾 �D�V�@@�@,�ЋD������Q�$�Q��h�  �R,�ҡD�������΋@�$h�  �@,�СD���jh�  �@�@0�СD���jh�  �@�@0�СD���jh�  �@�@4�и   ^]� U��V�uV�� �D�V�@@�@,�ЋD�����Q�$�Q��h�  �R,�ҡD���W��΋@�$h�  �@,�СD���j h�  �@�@4�СD�������΋@�$h�  �@,�СD���jh�  �@�@4�и   ^]� �������U��V�uV�C� �D�V�@@�@,�ЋD������Q��h�  h�  �R0�ҋD�jh�  �A�΋@4�и   ^]� �����U��V�uV�� �D�V�@@�@,�ЋD�W�Q���$h�  �Q�΋R,�ҡD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�и   ^]� ������������U��V�uV�� �D�V�@@�@,�ЋD�����Q�$�Q��h�  �R,�ҡD���j h�  �@�@4�и   ^]� U��V�uV胻 �D�V�@@�@,�ЋD������Q�$�Q��h�  �R,�ҡD������΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD���jh�  �@�@0�и   ^]� �������������U��V�uV�Ӻ �D�V�@@�@,�ЋD�W�Q���$h�  �Q�΋R,�ҡD���W��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD���j h�  �@�@0�СD���W��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD��@��j h�  �@0�СD�������΋@�$h�  �@,�и   ^]� ������������U��D�W�u�����   �O�@l�СD��u�O���   �@l�и   _]� ����U��V�uV�3� �D�V�@@�@,�ЋD���� �Q�$�Q��h�  �R,�ҡD���jh�  �@�@0�и   ^]� U��V�uV�Ӹ �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD�jh�  �A�΋@0�СD���j h�  �@�@0�СD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD���W��@�@,���$h�  �СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�и   ^]� ���������U��V�uV�� �D�V�@@�@,�ЋD�����Q�$�Q��h�  �R,�ҡD���j h�  �@�@4�СD���jh�  �@�@4�и   ^]� ����������U���V�uV耶 �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD�j h�  �A�΋@0�СD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@Qh<  �΋@8�СD��M�Q�@�@�Ѓ��   ^��]� ��U��]�g� �������U��V�uV�S� �D�V�@@�@,�ЋD������Q��jh�  �R0�ҋD�j h�  �A�΋@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���jh�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���jh>  �@�@0�и   ^]� ������������U���V�uV�� �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD�������A���$h�  �@,�СD��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M����@Qh<  �΋@8�СD��M�Q�@�@�Ѓ��   ^��]� �����������U��V�uWV�B� �D�V�@@�@,�ЋD�����Q�$�Q��h�  �R,�ҡD���W��ϋ@�$h�  �@,�СD���jh�  �@�@0��3����    �D���j �P��M  P�B4��F��|�D���jhY  �@�@4��_�   ^]� �U��V�uV胲 �D�V�@@�@,�ЋD�����Q�$�Q��h�  �R,�ҡD�������΋@�$h�  �@,�СD���j h�  �@�@4�и   ^]� ������������U���V�uV�� �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD�jh�  �A�΋@0�СD���j h�  �@�@0�СD���W��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD��M�W�fE�Q�E��΋@h�  �@H��(0�fE�D��M��p��E�Q�@��h�  �@H�СD��M�W�fE�Q�E��΋@h�  �@H�СD���jh�  �@�@0�и   ^��]� ������U���V�uV�`� �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD���W��A���$h�  �@,�СD�������΋@�$h�  �@,�СD���jh�  �@�@0�СD���jh�  �@�@4���� �E��tmj���� �E��t]�D�P�E�    �E��E�    ���   h�e P�A\�СD��M����@Qh�  �΋��   �СD��M�Q���   � �Ѓ��EP�Ċ ���   ^��]� �����U��V�uV�#� �D�V�@@�@,�ЋD������Q�$�Q��h�  �R,�ҡD���jh�  �@�@0�СD���jh�  �@�@4�и   ^]� ����������U��V�uV裮 �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD�jh�  �A�΋@4�СD���jh�  �@�@4�и   ^]� ��U��V�uV�3� �D�V�@@�@,�ЋD����X�Q�$�Q��h�  �R,�ҡD���� ��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD���jh�  �@�@0�СD���jh�  �@�@0�СD���jh�  �@�@4�и   ^]� �U���V�uV�`� �D�V�@@�@,�ЋD������Q��j h�  �R4�ҋD��A�M�Q�@�СD��M�j j�h���@Q�@�СD��M����@Qh<  �΋@8�СD��M�Q�@�@�Ѓ��   ^��]� ���������������U���u赬 �D��u�@@�@,�ЋD����ЋA��jh>  �@0�и   ]� U��V�uV�s� �D�V�@@�@,�ЋD������Q��j h�  �R0�ҋD�j h�  �A�΋@0�СD���W��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD���W��΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD�������΋@�$h�  �@,�СD��@������@,���$h�  �и   ^]� ���������������������������U��V�uV�� �D�V�@@�@,�ЋD������Q��j h�  �R0�ҋD�jh�  �A�΋@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���jh�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h�  �@�@0�СD���j h/  �@�@0�СD���j h0  �@�@0�СD���jh  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j hG  �@�@0�СD�j hH  �@�@0���СD���j hI  �@�@0�СD���j h  �@�@0�СD���j hK  �@�@0�СD���j hL  �@�@0�СD���j hM  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD��@��j h%  �@0�СD���j h&  �@�@0�СD���j h3  �@�@0�СD���j h4  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h'  �@�@0�СD���j h(  �@�@0�СD���j h5  �@�@0�СD���j h6  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h)  �@�@0�СD���j h*  �@�@0�СD���j h7  �@�@0�СD���j h8  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD���j h  �@�@0�СD��@�@0��j h  �СD���j h+  �@�@0�СD���j h,  �@�@0�СD���j h9  �@�@0�СD���j h:  �@�@0�СD���j h  �@�@0�СD���j h   �@�@0�СD���j h!  �@�@0�СD���j h"  �@�@0�СD���j h-  �@�@0�СD���j h.  �@�@0�СD���j h;  �@�@0�СD���j h<  �@�@0�СD���jh  �@�@0�СD���j hA  �@�@0�СD���j hB  �@�@0�СD���j hC  �@�@0�СD���j h  �@�@0�СD���j h1  �@�@0�СD���j h#  �@�@0�СD���j hD  �@�@0�СD���j hE  �@�@0�СD���j hF  �@�@0�СD�j �@�@0��h$  �СD���j h2  �@�@0�СD���j h  �@�@0�СD���j h
  �@�@0�СD���j hJ  �@�@0�СD���j h=  �@�@0�СD���j h>  �@�@0�СD���j h?  �@�@0�СD���j h@  �@�@0�СD���jh>  �@�@0�и   ^]� ��������������U���0V��E��MP�oF(ǆ�      ���   �E��oF8�E��w� �oM�W��o ǆ�      ǆ�       ���   ǆ�       f(�ǆ�   �����\U��\��M�\��E�\�f����   ^��]� ����������A    �   �A    �������������V���F\    ǆ�       �FX    ������vP�N �FT�R���   ^�������������A8���$��  �   ���������U���V���2@ ��u^��]ÍM��	 �D��M�htxt heman�@�@4�ЍE�Pj�N�9G h�  ���mC �M��5	 �   ^��]������������U���8V��~P ��   �FHW��oN(�E�M�E��oF8P��  �E؉�  �E�f(�  �\V0�\���  QP�N ǆ      �U��E�������@�YM�ǆ      �YE��XM��XE�f��oE��  ��(  ^��]� �������������U��E�A �EH��wb�$�غ�A$    �=�A$   �4�A$    �+�A$0   �"�A$@   ��A$P   ��A$`   ��A$p   �A0   �A,   �A(    �E�A   �A]� �I i�r�{�������������������U���0�D�S�]V�@��Wj hvdpi���   ���ЋD���j hacpi�Q�ˋ��   �҉E��E�    �E    ��suom�S  hTCAb�M��� �M��� ���T1 �D�Phdiem�Q�M�B4�СD��M�j havem�@�@4�Ѓ}���  �D���j hxvpi�@���   �ЉE��ˡD�j hyvpi�@���   �ЉE�΍EP�E�P�59 j ���F   ��/ �F ��t�u�u�jV�v�Ѓ��EЋ�Pjhsuom�[1 ����   �I �D��M�j havpi�@���   �Ѕ���   �D��M�j hxvpi�@���   �ЉE��MСD�j hyvpi�@���   �ЉE�΍EP�E�P�8 j ���L/ �F ��t�u�u�jV�v�Ѓ��D��M�jhrdem�@�@4�ЍE��P�/ �EЋ�Pjhsuom�0 ���8����D��M�j hrdem�@�@4�ЍE��P�v/ j ���F    ��. �F ��t�u�u�jV�v�Ѓ��u����u��P,��t2�~ t3�9F���Fj ���. �F ��t�u�u�jV�v�Ѓ��M�� �M��� _^�   [��]� _^3�[��]� ��U��D�V�uW�@��j hvdpi�΋��   ��=byekuV���.���_^]� =suomu6�D���j hbdpi�@���   �Ћ�V��t�����_^]� �a���_^]� _3�^]� ���U��Q���E��xP u3���]� S�]��u	3�[��]� W�}��j�k� ��t
_3�[��]� Vj��胘 �D�j W�@@�@8�Ѓ��E3����V�R\��t.V���7� ��t"V���+� ;�t!V���� �M�PS�e�����uF��c}�E�^_�   [��]� ^_3�[��]� �������������V��  �t?��   t6�����  c��u��  ��  �����^���  ��  �����^�3�^��U��� SVW���0� �Ѕ�t8�D�h-� R�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E���E�    �����aA ��3���~V���A F;�|���9 �E�3��E��E�    �H����   �D����   �@X�Ћ���t|��$    �M��( ���!� �D�Pheman�Q�M��B8�СD��M�Wheert�@�@p�ЍE���PV�h@ ���� ��t�M�V�$6 �u��誶 �M���F� ��u��u����!A ���J> j �u���A �E�P�9 ��_^[��]������������U��D��M����@VW�u�@(Q�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]����U��QSW���G    �l� �؅���   �D�h-� S�JL���   �ыЃ�����   �D�Vj R�A@�@8�Ћ������~   ���(����E���tpP���y�������tb�I � uHVS��������t+�D��΋��   �@�СD���j h�� ���   �@���u����� ����u�j j h,� �� ��^_[��]�����������U���DSVW�}����  �D�h-� W�@L���   �ЋЃ�����  �D�j R�A@�@8�Ћ؃��]����  �u����  �D�h-� V�AL���   �ЋЃ����z  �D�j R�A@�@8�Ѓ��E����[  � �E����2  �D�WP�I|�A$�Ѓ����  ���� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�ЋK�����:  �D����   �@X�Ћ؅��   �d$ �D����u�j ���   � �ЋM�jP�E���
 j �u��j,�>� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�ЋM��S�F���������  �D����u�j ���   � ���u�ȉE��ُ �D��E��u����   �H�Rh�ҋMj �u�j,�� �D��M�Q�@�@�СD��M�j j�h ��@Q�@�СD��M�Q�@�@�СD����΋��   �@��-�� t	��&��   �D�V�@@�@,�Ѓ���Wh�  �� �Ѕ���   �D��u�j ���   �ʋ �ЋM��j j W�a� �Mj Wj,��� �D��M�Q�@�@�СD��M�j j�h,��@Q�@�СD��M�Q�@�@�СD��u��@@�@,�ЋD����ЋA��Wh�  �@p�Ћ}S��肇 �����|�������� �u�؅�������D�j�u��@|�@,�Ѓ����� �D��M�Q�@�@�СD��M�j j�h8��@Q�@�СD��M�Q�@�@��j ��� j j h�� �� ��(�E��   P�� ����_^[��]� �E�3�P�� ����_^[��]� _^3�[��]� ����U��D����@SVW�}��@ ���Ћ]=fnic�  �~X ��   �~P �t  �D���j j�@���   �ЉE�ϡD�j j�@���   �ЉE�΍EP�EP��. fnM��fnE���j �������f���E�P�4  ���   P�E�P�$�������t�oE�E��j ���   ���   ��$ �}� u�E��t	����  �D���hfnic�@�@$�СD���jj�@�@4��SW����" _^[��]� �D��ϋ@�@ ��='  �g  �D���j j�@���   �Ѕ��I  �E��ΉE�EP�E�PW�. �}��   �  �M���  �D�j�hG  ���   ���   �Ѕ�u%�D��Mj�h�� ���   ���   �Ѕ���   j���. �D���j j�@���   �Ѕ���   �M�����3��E��E    ���~   ���D�W���   �M���   �ЋD��؋��   �ˋR��=G  t�D����   �ˋ@��=�� u�~P u���u�����t�u��S�v.���Ej ���J# G;}�|��   _^[��]� j����- SW���4! _^[��]� �����������U����}S��u=�M�E�Pj �E��  �E�    �E�    �~U ���GQ ��tj h&� �� ���u���u�u� [��]� �������������U��Q�}���E���   �D�V�u�@@�@,�ЋD�W�Q���$h�  �Q�΋��   �������W��\$�$h�  V�K& �D�������΋@�D$W��$h�  ���   ��������$h�  V�& �E���^�u���u�u�?� ��]� ���������U���SVW�}�ك���   ��Ҵ ��  �H� �D����u�I@�I,�у��E�V��h�  ����� ����  ��  �I �D���j W�@���   �Ћ3PW�r6������P�Vp�u�G���  ~��B  ��� �ȉE��� �D��E�P�I�I�ѡD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��u�@@�@,�ЋM�����u��	j �hS �8��0�����w*�D���j W�@���   �Ћ3PW�5������P�Vp�u����  uL�u���W�� ��t=��  ��I �D���j W�@���   �Ћ3PW�r5������P�Vp�u�G���  ~͋M���� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��u���u�u�F� _^[��]� �������������U��E��S�]V��W����   =Ҵ �L  �F� �D���S�I@�I,�у��؋ˉ]�Wh�  ��� ���  ��  �I �D���j W�@���   �Ћ��PW�RpG���  ~ٻ  �d$ S�J8���D������Q�M�j W���   �ҋ��PW�RpC��M  ~��  �� �ȉE��x� �D��E�P�I�I�ѡD��M�j j�h8��@Q�@�СD��M�Q�@�@�СD�S�@@�@,�Ћ؃��E�]�j ��9Q �8�}���0�����w �D���j W�@���   �Ћ��PW�Rp�8��������Iw-W�h7���D������Q��j W���   �ҋ��PW�Rp�}����  u}�u���W�^� ��tn��  ��I �D���j W�@���   �Ћ��PW�RpG���  ~ٻ  �d$ S��6���D������Q�M�j W���   �ҋ��PW�RpC��M  ~̋M��D� �D��M�Q�@�@�СD��M�j j�hH��@Q�@�СD��M�Q�@�@�Ѓ��E�]�u��PS賎 _^[��]� ����������U��D����@V�uW�@ ������=TCAb��   �D���j hdiem�@���   ��=�  ��   �D���j hghcv�@���   �Ѕ�u=�D�������΋@�$havem���   ���]��E�f.�����D{>�D���W��΋@�$havem���   �Ѓ����]��E��G8�$�m�  �u��V�f _^��]� ����������U��]��) �������U���<  SVW���P ��  �� �ȅ�t7�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3��oEj ���ϋ�� �E�P�  j�wP����5���oE�E���   H��  Ht#H�f  9E$�]  j�� ��_^[��]�$ �}$ tAj��������P�{��j ���o ������P���   �~{���o ���   _^[��]�$ �} ��  �}  ��  �E�H����  �$����M�����  jj j��� �M��#� j h���M������D��M�Qh�� �M�@�@8�СD��M�Q�@�@�Ѓ��M�j h��������D��M�Qh�� �M�@�@8�СD��M�Q�@�@�Ѓ���D���j h�������D���D���Qh�� �M�@�@8�СD���D���Q�@�@�Ѓ���T���j h���T����D���T���Qh�� �M�@�@8�СD���T���Q�@�@�Ѓ���$���j h������P��t���蓿���D���t���Qj �M�@���   �СD���t���Q���   � �СD���$���Q�@�@�Ѓ��M�j h��諿���D��M�Qhô �M�@�@8�СD��M�Q�@�@�Ѓ���4���j h���l���P�M������D��M�Qj �M�@���   �СD��M�Q���   � �СD���4���Q�@�@�Ѓ���d���j h�������D��@��d���Qhɴ �M�@8�СD���d���Q�@�@�ЋG�M�j j
Qh���h����p�af ����~j j P��� ���M��� _^[��]�$ �u����+  j �wP���u2��jj j���H j �/j j�j �+�u�����  j �wP���E2��jj j��� �u��u�Vh���h������`�  _^[��]�$ �}$ �Z����} �E���   H��   HtQH��  �u�����  �}�c��  j �E$�E$����PV���U�  �؅���  �u$��jj V�~ VS��  �u����D  j �wP���1��jj j���a~ V���ɨ  �(  �}  t;HtUH�  �u����  P���qy ��jj ����   j �~ _^[��]�$ H����  �$���j �wP���1��E�G\   E��oE��G`�Gp_^[��]�$ �}� tmj�R� �D������   ���   �Ћu���j �E$��x ��tj �u$�Ϟ�����	�M$V�A���j �u$��h�   �u(��  �M$�����_^[��]�$ �u����  j ���x ��uP�wP���Y0��jj ��j�,} �oE���ϋ�V� �����_^[��]�$ �}� ��  �u�����  �E�E$�����  �OP�!� �]��M�f.�����DzW�fE��E��E��E��E���E�^��E��E�^��EԋOP�����P�R� �E̋��X �E��@�������XE�P�E���x �E̋M��\ �E��E��\@������P�E��x �]��U��M��\P�\�E��Y��Y��Y��Y��X��X�f/�v�u��c   �E$��E��t=��cu8j�`� ������jcV�oE���ϋ�� � ���_^[��]�$ �]�u���]$j�%� ����tX��ct�S���av �E$��tjj S����z jc�u$�S랋M������j@P�z P�]� �D������Q�@�@�Ѓ�_^[��]�$ ����������A�i���������U���(V��VP����  �M��HtH�  H�~  �}$ ��  �FH�E�P���E�臟 �]�\��   �F`�U�\��   fW`��\�fW`��F`�Fh�\��Fh�Fp�\��Fp�Fx�\��Fx��  �\���  ��   �\���   ��(  �\���(  ��0  �\���0  �E�f.�����D��   W�fE��U��]���   �}$ �u  j �E��P��r���E����\��   �$�VC���]��M���fW`�f.�����D�)  �o��   �����vP� ���$�Po �]��E��N �Y ��XFH�$�η  �oE����   �oE���   ^��]�  �^��^��M؃��E��XˋNP�X�f���^� �oE���   ^��]�  ��u}�~\ t'�oEj ���Fp蜣  �oE���   ^��]�  ���    t)�oE���΋�� �J/���oE���   ^��]�  ��    t�oE���΋�� ����oE���   ^��]�  ����U���SV��W�~P ��  �� �؅�t7�D�h-� S�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3��EHtGHt$H��  9E$��  PPhƴ �2� ����  �} ��  j j hǴ �� ���  �~\ t	j���k�  ��    t(��   t��  ����  ��  ��  �:������   �Z  ���� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ���j ���   j*�� �D��M�Q�@�@�СD��M�j j�h ��@Q�@�СD��M�Q�@�@�Ћ��   ��j���   j �"v j ���   ��j*�A� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ћ��   ��j���   ���   �u ����� �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ѓ�j�vP���F\    ǆ�       ǆ       ǆ�      ��(��j�K� �D����   ���   ��j P�E�ݖ���u�M����= Pj Vh+� �Qf ���M��&@ �D��MQ���   ���   �Ѓ�_^[��]�  ���U����} VW��tL�}  �
   �NP�   E��E�P�� ����} fn����}�M��\��M��\�XE��E��P�}$ th�}  �
   �NP�   E��E�P衙 ����} fn����}�M��\��M��
�XE��E��oE��NP����� ��� _^��]�  �E��yj j hŴ �~j j hĴ ��� ��_�FX    �F\    ǆ�       ǆ       ǆ�      ^��]�  �������������3���������������U����   �D�V��W�@j �FH�NT���   �E��oF(hT  �u���H����oF8��X����Ћ��K� �ȅ�t7�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3�WɍGf(��}�\�H����vP�   �G    �E��E�f(��\�P���fn�����G�����G    �G    �E��YM��E�f(��M�fW`��E�f(��Y��E��y}�����u؅��n  E�E�d$ �D�j V�@@�@8�ЋM����E��x���VP�I �w�����x���������Y����P�E��E��Y���E���n �E���x����U�� �\e��X�\]��m�M�Y��Y��Y��Xe��X]��Y��E�� ����E�f/��u��e��]���$����k  (��X�f/���8����R  �� ���f/��@  �X�f/���(����*  �M���h���VP�I �o�����h�����X����Y����P��@�����p����Y����0�����m �M���h�����p���� �X�\�@����\�0����AH�i(�Y��Y��Y��Y��A8�X�f/���   �X�f/�wv�Q0�A@�X�f/�wb�X�f/�wX�M�m�]��E�e�f/��E��e�r,��8���f/�v�U��M�f/�r��(���f/�wU�E����pP��j ���E؅�������?�N  �E�W��M�U�\M��\U�f.ß��D�u  W��  �E��}��X��XM�f(��   �w�e��X��M��]��M��M��E��E��U���E�X��f(��M�X���E�f/�r5�E��X�f/�v&�M�f/�r�X�f/�v�G   ��_^��]� �E܋�P�-n �D��ЋA�ʋ@<�ЋD�����E�P�I�I�у�����   �E��XE��e��E��E��U��E��E��]��M���E�X��U���M�X��]�E��E�f/��E�r4�E��X�f/�v%�M�f/�r�X�f/�v�   ��_^��]� �M��@T�Ѕ���   �M���X���jc�u�P�I �!����e�� �YE��H�YM��XE��XM��E��U��E���E�X��U��M��]��M���M�X��]�E��E�f/��E�r;�E��X�f/�v,�M�f/�r!�X�f/�v�   ���Gc   _^��]� �M3���@d�Ѕ��J����MV��@\�Ѕ���   �M���X���V�u�P�I �/����e�� �YE��H�YM��XE��XM��E��U��E���E�X��U��M��]��M���M�X��]�E��E�f/��E�r$�M��X�f/�v�E�f/�r
�X�f/�w�MF��@d��;��&����k����   �ǉw_^��]� �^��^��M��U�fE܋u���j ����� ��T���P�����o �@��G�?ui�U�W��E�M�\E��\M�f.ӟ��DzW���^��^��E��M�fE�j ���΋�� ��T���P������o �@��G��_^��]� �������������U����   SV��W�u��z� ���}���t:�D�h-� W�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E����3ۉ]��]� �E�D����   ���   �ЉE��E����  �D�WP�I|�A$�Ѓ�����  �u������C���M��E��D����   ���   �Ѕ���  ��蘻 �D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�Ѓ���j �vP�����D�W��NTj hR  �@fE����   �ЋD��؋NTj hZ  �R�]����   �҉E����Y  �D�3�(@��M�fE싀�   (p�fE����   ���U����   �E��E��E��E��E��U��EȡD��M�V���   ���   �ЍM�Q���f �M��E�f/�v�M��E��U�f/�v�E�f/M�v�M�f/E�v�EСD�F�M����   ���   ��;�|��E��M��U��]���]��E��M��\u��\��Y���Y���X��X��E��M��E��E��E��E��E��E��E��E��D�3ۋM��]̋��   ���   �Ѕ��  �I �D��M�S���   ���   ��j �؋�Sj(蛹 �D��A��8���Q�@�СD���8���j j�h��@Q�@�СD���8���Q�@�@�СD����ˋ��   �@L�СD��M�S���   �@h��j Sj,��� � �D���X���Q�@�@�СD���X���j j�h��@Q�@�СD���X���Q�@�@�Ѓ����vP��h jj j���h �E�P���d �E���u&�M���E���\M��\E�f����   ��uv�NP��(���P赍 �NP� �Y���E��@������Y��P�E��c� �U��]��M��@�\U��X�XE��\M��X��X�f��B��uMj��x�����P�y`���E��\E��M��\M���x����X��E��X�fЃ�������lh �vP���2b �D�������IV�I�ыD�VW�A�@�ЋM��E���P�}�  �}���j Sj(�n� �D���H���Q�@�@�СD���H���j j�h(��@Q�@�СD���H���Q�@�@�Ѓ��E���P�Kf �D�S�@@�@,�ЋD����EԋQ��jh�  �R0�҃}� �  �D��ˋ��   �@��-�� t	��&��   �D��ˋ��   �@��=�� uhG  �"�D��ˋ��   �@��=մ ��   h�� �m� ��������   j j V���ԡ j Vj,���X� �D���h���Q�@�@�СD���h���j j�h4��@Q�@�СD���h���Q�@�@�СD����Mԋ@Vh�  �@p�СD���j hҴ ���   �@�СD��M�Q�@�@�СD����]̋M�C�]̋��   ���   �Ћu�;�������D�j�u�@|�@,�ЋM��W��������`� �D��M�Q�@�@�СD��M�j j�h@��@Q�@�СD��M�Q�@�@�Ѓ��J�D��M�Q�@�@�СD��M�j j�h���@Q�@�ЍE�j P�i� �D��M�Q�@�@�Ѓ� �D��M�Q���   ���   �ЍE��E�    P��� ��_^[��]�����U��E��
wQ�$�d�3�]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø   ]ø	   ]ø   ]Ã��]ÍI ���$�+�2�9�@�G�N�U�U��E��
wT�$�����  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]ø�  ]Ã��]â���������������������U��E��H�  �$�<��/  ]ø0  ]ø  ]ø  ]ø  ]øG  ]øH  ]øI  ]ø  ]øK  ]øL  ]øM  ]ø  ]ø  ]ø  ]ø  ]ø  ]ø  ]ø%  ]ø&  ]ø3  ]ø4  ]ø  ]ø  ]ø  ]ø  ]ø'  ]ø(  ]ø5  ]ø6  ]ø  ]ø  ]ø  ]ø  ]ø)  ]ø*  ]ø7  ]ø8  ]ø  ]ø  ]ø  ]ø  ]ø+  ]ø,  ]ø9  ]ø:  ]ø  ]ø   ]ø!  ]ø"  ]ø-  ]ø.  ]ø;  ]ø<  ]ø  ]øA  ]øB  ]øC  ]ø  ]ø1  ]ø#  ]øD  ]øE  ]øF  ]ø$  ]ø2  ]ø  ]ø
  ]øJ  ]ø=  ]ø>  ]ø?  ]ø@  ]Ã��]Ë�6�=�D�K�R�Y�`�g�n�u�|������������������������������������������$�+�2�9�@�G�N�U�\�c�j�q�x������������������������������������������ �'�.�U��W��j�u�O�-� �Oj�u� � �   _]� ������U���TVWh+  �> �D����E�P�I�I�ыD��A�M�QV�@��jh��jxj�Ǧ ���� ��t���� ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P��� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �Z �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��	� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh	+  �. �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j贤 ���� ��t���Ԣ ���3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P��� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Phɴ �G �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M���� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���TVWh�*  � �D����E�P�I�I�ыD��A�M�QV�@��jh��jj觢 ���� ��t���Ǡ ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �: �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M���� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh�*  � �D����E�P�I�I�ыD��A�M�QV�@��jh��jj藠 ���� ��t��跞 �l��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �*� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M���� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh�*  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��j0j臞 ���� ��t��觜 �@��3��D��M�Q�@�@�СD��M�j j�hd��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M���� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh�*  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��jHj�w� ���� ��t��藚 ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �
� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh+  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��jTj�g� ���� ��t��臘 ����3��D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�x� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Phô ��� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh +  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��j`j�W� ���� ��t���w� � ��3��D��M�Q�@�@�СD��M�j j�hD��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�h� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh�*  �  �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j�D� ���� ��t���d� ���3��D��M�Q�@�@�СD��M�j j�h(��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�U� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���TVWh�*  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��j$j�7� ���� ��t���W� ���3��D��M�Q�@�@�СD��M�j j�h0��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�H� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� ��� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��y� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh+  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��jlj�'� ���� ��t���G� �\��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�8� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��i� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]�����������U���TVWh+  �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j�� ���� ��t���4� ����3��D��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�%� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�PhǴ �� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��V� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���TVWh�*  �~� �D����E�P�I�I�ыD��A�M�QV�@��jh��j<j�� ���� ��t���'� �t��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph�� �� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��I� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]���������������������������U���TVWh+  �^� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j�� ���� ��t���� ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P��� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Ph´ �w� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��&� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���TVWh+  �N� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j�ԉ ���� ��t���� ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�� �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�Phƴ �g� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���TVWh+  �>� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j�ć ���� ��t���� �<��3��D��M�Q�@�@�СD��M�j j�h`��@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�պ �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�PhĴ �W� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M��� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���TVWh+  �.� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j贅 ���� ��t���ԃ �p��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ�(�E��M�P�Ÿ �M�Q�0�D��@�@�СD��M�Q�M�Q�@�@�СD��M܃��@�@<�ЋD�j�j��Q�MQP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�Ѓ��D��M�@�@<�ЋD�j�j��Q�M�QP�M�BL��W�E�PVj �E�PhŴ �G� �D����E�P�I�I�ыD��A�M�Q�@�Ѓ� �M���� �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��MQ�@�@�Ѓ���_^��]��������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��hR  j襃 ���� ��t���Ł ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phl� �� ���M����޶ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��hs  j�e� ���� ��t��� �D��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hh��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M�襳 V�M�Q�0�E�h   Pho� ��� ���M���螴 �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h  j�% ���� ��t���E} �D��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hh��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��e� V�M�Q�0�E�h   Phf� �� ���M����^� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh̴ �_� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j��| ���� ��t���{ ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��%� V�M�Q�0�E�h   Phy� �K� ���M����� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h  j�z ���� ��t����x �|��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phg� �� ���M����ޭ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhT� ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��h{  j�ex ���� ��t���v ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M�襪 V�M�Q�0�E�h   Ph�� ��� ���M���螫 �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h]  j�%v ���� ��t���Et ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��e� V�M�Q�0�E�h   Phm� �� ���M����^� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �_� �D����E�P�I�I�ыD��A�M�QV�@��jh��h&  j��s ���� ��t���r ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��%� V�M�Q�0�E�h   Phh� �K� ���M����� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhN� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��hO  j�q ���� ��t����o ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h ��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Ph�� �� ���M����ޤ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��h~  j�eo ���� ��t���m �|��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M�襡 V�M�Q�0�E�h   Php� ��� ���M���螢 �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhִ �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h.  j�%m ���� ��t���Ek �,��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hP��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��e� V�M�Q�0�E�h   Ph�� �� ���M����^� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �_� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j��j ���� ��t���i ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��%� V�M�Q�0�E�h   Phq� �K� ���M����� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�h ���� ��t����f ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phr� �� ���M����ޛ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�ef ���� ��t���d �4��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hX��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M�襘 V�M�Q�0�E�h   Phs� ��� ���M���螙 �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhʴ �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h1  j�%d ���� ��t���Eb ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��e� V�M�Q�0�E�h   Phi� �� ���M����^� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhO� �_� �D����E�P�I�I�ыD��A�M�QV�@��jh��hZ  j��a ���� ��t���` ���3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h<��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��%� V�M�Q�0�E�h   Ph�� �K� ���M����� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h<  j�_ ���� ��t����] �(��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hL��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Phj� �� ���M����ޒ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhϴ ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�e] ���� ��t���[ ���3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h(��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M�襏 V�M�Q�0�E�h   Ph{� �˻ ���M���螐 �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]������������������������������U���dVhʹ �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�[ ���� ��t���5Y ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��U� V�M�Q�0�E�h   Phz� �{� ���M����N� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhS� �O� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j��X ���� ��t����V �<��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h`��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Ph�� �;� ���M����� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhѴ �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h  j�V ���� ��t���T �x��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��Ո V�M�Q�0�E�h   Ph}� ��� ���M����Ή �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �Ͼ �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�UT ���� ��t���uR �T��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hx��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M�蕆 V�M�Q�0�E�h   Phx� 軲 ���M���莇 �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� 菼 �D����E�P�I�I�ыD��A�M�QV�@��jh��hG  j�R ���� ��t���5P �`��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��U� V�M�Q�0�E�h   Phk� �{� ���M����N� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �O� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j��O ���� ��t����M �l��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Pht� �;� ���M����� �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhش �� �D����E�P�I�I�ыD��A�M�QV�@��jh��hD  j�M ���� ��t���K ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��� V�M�Q�0�E�h   Ph�� ��� ���M����΀ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �ϵ �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�UK ���� ��t���uI ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��} V�M�Q�0�E�h   Phu� 軩 ���M����~ �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� 菳 �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�I ���� ��t���5G ���3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h@��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��U{ V�M�Q�0�E�h   Phw� �{� ���M����N| �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhU� �O� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j��F ���� ��t����D � ��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h$��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��y V�M�Q�0�E�h   Ph�� �;� ���M����z �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh״ �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h9  j�D ���� ��t���B �h��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M���v V�M�Q�0�E�h   Ph�� ��� ���M�����w �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhQ� �Ϭ �D����E�P�I�I�ыD��A�M�QV�@��jh��hp  j�UB ���� ��t���u@ ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��t V�M�Q�0�E�h   Ph�� 軠 ���M����u �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� 菪 �D����E�P�I�I�ыD��A�M�QV�@��jh��hh  j�@ ���� ��t���5> ���3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h,��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��Ur V�M�Q�0�E�h   Phn� �{� ���M����Ns �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �O� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�   j��= ���� ��t����; ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��p V�M�Q�0�E�h   Phd� �;� ���M����q �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]������������������������������U���dVhԴ ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��h  j�; ���� ��t���9 ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M���m V�M�Q�0�E�h   Ph~� �� ���M����n �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhд 迣 �D����E�P�I�I�ыD��A�M�QV�@��jh��h  j�E9 ���� ��t���e7 �@��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hd��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��k V�M�Q�0�E�h   Ph|� 諗 ���M����~l �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� �� �D����E�P�I�I�ыD��A�M�QV�@��jh��h  j�7 ���� ��t���%5 ���3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h,��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��Ei V�M�Q�0�E�h   Phe� �k� ���M����>j �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhP� �?� �D����E�P�I�I�ыD��A�M�QV�@��jh��he  j��4 ���� ��t����2 �T��3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�hx��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��g V�M�Q�0�E�h   Ph�� �+� ���M�����g �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVh�� ��� �D����E�P�I�I�ыD��A�M�QV�@��jh��h�  j�2 ���� ��t���0 ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M���d V�M�Q�0�E�h   Phv� �� ���M����e �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U���dVhմ 迚 �D����E�P�I�I�ыD��A�M�QV�@��jh��h#  j�E0 ���� ��t���e. ����3��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�j j�h��@Q�@�СD��M�Q�@�@�СD��M܃�@�@Q�M�Q�@�СD��M܃��@�@<�ЋD�j�j��Q�M�QP�M܋BL�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�ЍE�P�M��b V�M�Q�0�E�h   Ph� 諎 ���M����~c �D��E�P�I�I�ѡD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���^��]��������������U��D��M��$�@VQ�@�СD��M�j j�h���@Q�@��jh��j:j�. ����$��t���., ����F    �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�Ca V�M�Q�0��h   Ph&� �j� ���M����=b �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�hx��@Q�@��jh��jEj�- ����$��t���>+ �T��F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�S` V�M�Q�0��h   Ph'� �z� ���M����Ma �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�h���@Q�@��jh��jPj�., ����$��t���N* ����F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�c_ V�M�Q�0��h   Ph(� 芋 ���M����]` �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�h���@Q�@��jh��j[j�>+ ����$��t���^) ����F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�s^ V�M�Q�0��h   Ph)� 蚊 ���M����m_ �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�h,��@Q�@��jh��jfj�N* ����$��t���n( ���F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�] V�M�Q�0��h   Ph*� 誉 ���M����}^ �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�hh��@Q�@��jh��jqj�^) ����$��t���~' �D��F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�\ V�M�Q�0��h   Ph+� 躈 ���M����] �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�h���@Q�@��jh��j|j�n( ����$��t���& ����F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�[ V�M�Q�0��h   Ph,� �ʇ ���M����\ �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]�U��D��M��$�@VQ�@�СD��M�j j�h���@Q�@��jh��h�   j�{' ����$��t���% ����F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�Z V�M�Q�0��h   Ph-� �׆ ���M����[ �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]��������������U��D��M��$�@VQ�@�СD��M�j j�h��@Q�@��jh��h�   j�{& ����$��t���$ ����F   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�Y V�M�Q�0��h   Ph.� �ׅ ���M����Z �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]��������������U��D��M��$�@VQ�@�СD��M�j j�hX��@Q�@��jh��h�   j�{% ����$��t���# �4��F	   �3��D��M�Q�@�@�СD��M�j j�h<��@Q�@�Ѓ��E܍M�P�X V�M�Q�0��h   Ph/� �ׄ ���M����Y �D��E�P�I�I�ѡD��M�Q�@�@�Ѓ���^��]��������������U���(S��W�]��3 �Ѕ�t5�D�h-� R�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��H��u3��}���D����   �@X�Ћ��E�3��E��E��A� ���E�P���#� ����   V��3�衊 ��~Q�3 �M؋��K �E؋�PV�R� �D�j Wheert�A�M؋@l�ЍM؋���K �E�;�to��F�P� ;�|��D��M�Q�@�@�СD��M�j j�h���@Q�@�ЍE�P�; �D��M�Q�@�@�ЋM���<H��^�E�P肂 ��_[��]Ë��  ��t5�D�V�u��@\�@,�Ѓ���u�M�� �M�V�% �E�   �u���u�M���  ���}���������E���t��D��M�Q�@�@�СD��M�Wj�h���@Q�@�ЍE�P�G: �D��M�Q�@�@�Ѓ����u��ɉ ���� WV���9� �E�^P证 ��_[��]�������U��SVW�}���u�|1 ���^����   �N0����   �D�Q�@�@�Ѓ�����   ���4�  ����   �D�S�@@�@,�ЋD����؋Q��j h�  ���   �҅�tm�D���j h�  �@�@0�ЋN0�[ �N0j jjZjZ�M\ �N0j j j �/] Wh�  ���bJ ��t j ���ER ��tj jh   �v0���\ _^[]� �������U���u��j h&� �;� ]� �������U��V�u��j h�� �� ����tj j h�� �&< ����^]� ������������U���V���W��f/��E��E��$v�G$ �� # �]��E�������FW�f/��E��E��$v�$ ���" �]��E����F���FW�f/��E��E��$v��# ��" �]��E����F���FW�f/��E��E��$v�# ��y" �]��E����F^��]�����U���@SVW���0/ �؅�t7�D�h-� S�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3�����( �D��M�Q�@�@�СD��M�j j�hT��@Q�@�СD��M�Q�@�@�ЋE��HK������  �$��|���̀���  j ����h���s  ����k���g  �������[  �vP����  �L  j �vP���֊���;  �������/  S�vP��芌���  �FH�E�jP���E����������o ��E��X ��1�FH�E�jP���E��{��������o ��E��\ ��vP�N ���$�  �   ���q ���+�����P��p �NP�+�����P��  j�E���P���������o �vP��N ������$�N  �F�vP����������t6�
��$    �I �D�j hȴ ���   �ϋ@���vP���<�  ����u֋���& �D��M�Q�@�@�СD��M�j j�h`��@Q�@�СD��M�Q�@�@�Ѓ���j �o _^[��]� ��{{'{3{�|?{N{_{�|�|�|k{{{�{|�{�|T|����U��W�}��t)VW��������tj j j����  W���c�  ����u�^_]� �������U��Q�D�SVW�@@�}j W�@8�M��Ѓ���3����V�R\��t'V���8�  ����tjj j���E�  �M�W�����}F��c|�_^[��]� ����������U���   W���P ��  �GHW��oW(S�E��oG8��h���f(��\O0�\��,��,؉E��]+ �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3�V�wP�������D����OTj h[  �R���   �҉E���L  �O V�E�P� ���E���h����Y����P�E��E��Y���E���  �U��u��_h��\M��@�\E��}��Y��Y��Y��u��M��Oxf/��E��Y�vf(��f(�f/�v�]���M��W`�Gpf/�vf(��f(�f/�v�U���E�f/�w(�f/�w(Ѓ}� �E��\e��\m�fn�����\�fn�����\��E�tO�X�f/��   �X�f/���   �E��X�f/���   �X�f/���   3�9Ej ��Pj��   �E��E��u��M��E��E��E��E��f/��E���   �X�f/�v{�E�f/�rp�X�f/�vf�E��XE��X}��E��u��M��}��E��E��E��f/��E�r&f/�v �E�f/�rf/�v3�9Ej ��Pj�jjj ���(�  �wP�����  ���O �������^[_��]� ��������U��IW�}��t4�D�V���   �@X�Ћ���t3���;���P��  �����  ����u�^�} tj Wh�� �4 ��_]� ���U����  �D��u�M�@@�@,�ЋM���E�j �� �8�  �P  �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��u���   �@8��H������  �$��j h�������4���D��M�Q�����Q�@�@�Ѝ�����  j h������������D��M�Q������Q�@�@�Ѝ������V  j h���M������D��M�Q�M�Q�@�@�ЍM��*  j h ���H�������D��M�Q��H���Q�@�@�Ѝ�H�����  j h��M��l���D��M�Q�M�Q�@�@�ЍM���  j h��������=���D��M�Q������Q�@�@�Ѝ������  j h(���h�������D��M�Q��h���Q�@�@�Ѝ�h����_  j h0���h��������D��M�Q��h���Q�@�@�Ѝ�h����*  j h8���H�������D��M�Q��H���Q�@�@�Ѝ�H�����  j hD��������i���D��M�Q������Q�@�@�Ѝ�������  j hT���(����4���D��M�Q��(���Q�@�@�Ѝ�(����  j hd���(��������D��M�Q��(���Q�@�@�Ѝ�(����V  j hl��M������D��M�Q�M�Q�@�@�ЍM��*  j hx�����������D��M�Q������Q�@�@�Ѝ�������  j h���M��l���D��M�Q�M�Q�@�@�ЍM���  j h���M��@���D��M�Q�M�Q�@�@�ЍM��  j h���M�����D��M�Q�M�Q�@�@�ЍM��q  j h����x��������D��M�Q��x���Q�@�@�Ѝ�x����<  j h����X�������D��M�Q��X���Q�@�@�Ѝ�X����  j hļ��8����{���D��M�Q��8���Q�@�@�Ѝ�8�����  j hм������F���D��M�Q�����Q�@�@�Ѝ�����  j hܼ����������D��M�Q������Q�@�@�Ѝ������h  j h������������D��M�Q������Q�@�@�Ѝ������3  j h�����������D��M�Q������Q�@�@�Ѝ�������   j h���������r���D��M�Q������Q�@�@�Ѝ�������   j h����x����=���D��M�Q��x���Q�@�@�Ѝ�x����   j h���X�������D��M�Q��X���Q�@�@�Ѝ�X����bj h���8�����
���D��M�Q��8���Q�@�@�Ѝ�8����0j h �������
���D��M�Q�����Q�@�@�Ѝ�����D�Q�@�@�Ѓ��D��M�Q�M�h<  �@�@8�СD��M�Q�@�@�Ѓ��u�M��u�u�u���  ��]� ����/�d���ł�&�[���Ń��/�d���ń��I�~�����R������&�X�����������U���X�D�SVW�@@�u�M��@,�Ћ]�����ˉ}�j ��� �8�  �z  �D��u���   �@8�ЋD������Q��j h�  ���   �ҋD����E�P�I�I�ыD�j j�h��A�M�Q�@�ЋM��E���VP�#����D����E�P�I�I�ыD��A�M�QV�@�СD��M؃��@�@<�ЋD�j�j��Q�M�QP�M؋BL�ЋM��E�WP������D����E�P�I�I�ыD��A�M�@Q�M�Q�СD��M���@�@<�ЋD�j�j�V�Q�M�P�BL�СD��M�Q�M�h<  �@�@8�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�ЍM���   j ���Q� �8�  �	  �D���j h�  �@���   �ЋD����u���   �I8�ыD����E�P�I�I�ыD�j j�h��A�M�Q�@�ЋM��E��VP藿���M�P�E�PW�E�P腿��P�E�P�����P�E�P�����D����Q�M�Ph<  �B8�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�ЍM�D�Q�@�@�СD��M�Q�@�@�Ѓ��u�M��uS�u�Z�  _^[��]� �U���   �D��u�M�@@�@,�ЋM���E�j ��� �8�  ��  �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��u���   �@8�Ѓ����  �$�ȍj h|���x����%���D��M�Q��x���Q�@�@�Ѝ�x����2  j h���M������D��M�Q�M�Q�@�@�ЍM��  j h���M������D��M�Q�M�Q�@�@�ЍM���   j h���M�����D��M�Q�M�Q�@�@�ЍM��   j h���M��o���D��M�Q�M�Q�@�@�ЍM��   j h���M��C���D��M�Q�M�Q�@�@�ЍM��Yj h���M�����D��M�Q�M�Q�@�@�ЍM��0j h����h��������D��M�Q��h���Q�@�@�Ѝ�h����D�Q�@�@�Ѓ��D��M�Q�M�h<  �@�@8�СD��M�Q�@�@�Ѓ��u�M��u�u�u��  ��]� 	�>�j�����@���������U���x�D��u�M��@@�@,�ЋM���E�j 臐 �8�  ��  �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��u���   �@8�Ѓ����  �$�ȏj h��M�����D��M�Q�M�Q�@�@�ЍM���   j hм�M�����D��M�Q�M�Q�@�@�ЍM��   j h���M��c���D��M�Q�M�Q�@�@�ЍM��yj hܼ�M��:���D��M�Q�M�Q�@�@�ЍM��Pj h��M�����D��M�Q�M�Q�@�@�ЍM��'j h��M������D��M�Q�M�Q�@�@�ЍM��D�Q�@�@�Ѓ��D��M�Q�M�h<  �@�@8�СD��M�Q�@�@�Ѓ��u�M��u�u�u��  ��]� v���Ύ�� �I�U���H�D�V�u�M��@@�@,�ЋM���E�j 薎 �u�8�  �,  �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD�V���   �@8�ЋD�P�E�P�I�A(�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M��<�@�@<�ЋD�j�j��Q�M�QP�M�BL�СD��M�Q�@�M��@8h<  �СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ћu���u�M�V�u�u�y�  ^��]� ��U��D�V�uW���   ���FP�B<��3����_8�>���G@�   _^]� ������U���h���@�Mf/�VW��w��f/�v(�(��^F(f.���E���D�T  �}�E�P���N(���  �E���P���  �m�W��M��E��u�}f(��\]��f(��\U�f.��E��E��E�W��fE���D{	�^��]��E�f.ğ��D{	�^��U��Ef.ğ��DzW�fE��U��]���]��U��^��^��m��M��E��f.��E��E��E��E���Dzf.ğ��DzW�fE��U��]���Y��Y��\���\��ċ�f��0�[�  �F(�����$��  W����,��_^��]� �������U��S�]V��9^P��   W�7 �ȅ�t7�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ����3�S�N �^P�|,���FP��t1jP���K���j j hɴ �! j �vPh�� �! ��_^[]� j j h�� �! ��_^[]� ������������U���P�D�W�VW�����@�$�O ���   j	�СD��O ��W��]��@�$j���   �СD��O ��W��]؋@�$j���   �СD��O j j�]�@���   ��j j���E��  W��E�    ���ύE�$V�E��� �D$�E��D$�E��D$�E�$P�j �D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ���rgdft{��tcpf��   �D��M��E�Yp�Q�@�E�@�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�ЍM��u�E�M��Y���D�Q�^(��@�@�E�СD��M�j j�h���@Q�@�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�ЍM�D�Q�@�@�Ѓ��D��M��Ej0j �@j	j����@$�$Q�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@���E��,W�f.����D�D��@zQ�@�M�Q�СD��M�j j�h���@Q�@�СD��M�Q�M�Q�@�@�СD��M�Q�@�@�Ѓ� ��   �@<�M��Ѝp���~!�D�V�A�M�Q�@4�Ѓ�f��0uN��ߡD��M�VQ�@�@4�Ѓ�f��.uN�D��M��P�FPj �E�P�BP�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M�Q�@�@�Ѓ��D��M��E�  �E    Q�@�@�СD��M�Q�M�Q�@�@�СD��MЃ��@�@<�ЋD�j�j��Q�M�QP�MЋBL��j j �EЋ�P�EP�l �D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ�_^��]� ��U���TSVW���}�� �ȉM���t8�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E���E�    �D����j j �@�@�Ћ؋�j�E��]�P�L����} �.  �D�3�������   �@X�ЋЅ��  �D�F���   �ʋ@(�ЋЅ�u����   �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M��E�    �E�    Q���   �M�Q�@$�СD��M����@Qj �ˋ��   �СD��M�Q���   � �СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��MЃ��@Qh�� �ˋ@8�СD��M�Q�@�@�Ѓ��Gj j
S�u�u�p螟 �u���؉]��t���H( V��  ������  �D��M�Q�@�@�СD��M����@QS�M����   Q����ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M�Q�@�@�СD�������P��'  j P���   �Ѓ} �Euj�E���P�#����o ��oE��M��E��K �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�Ѓ��M���& �E�Phacpihbyek�!� �D��M����@j haqpi���   �ЍM�����& ��u�M�V�����M�P�cj���E3�=�� uSSP� ���/  =�	 ��   �oE������u�� �D�jj ���@��V�@�СD��M�VQ�@�@�ЋM���h�� �r  �؅���   �D�S�@@�@,�ЋM��Q�� �D��������   ��j V���   �ҋD�Vh�  �A�ϋ@p�СD�j S�@@�@8�Ѓ��ȋj �Rh�e�M��-�� t+��&t����Q�:h�� ���8W���؅�u:����hմ �hG  ���W���؅�u����h�� �oE���� �Y���؋u����   ���~   �D�j S�@@�@8�Ѓ����} t.���j �R\��tj�u��j �/�  ����PT��t=jS�u�.�E��cu"3������V�P\��uF��c|��j�u��V�jSP����  �M�j �MN �M��� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M�Q�@�@�СD��M�Q�@�@�ЋE��_^[��]� _^��[��]� ��������������U���@VW�M��` ���M��u���# ��u�M�����D$ ��_^��]� �D�Sh-� V�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��E����3ۉ]��K��u3���D����   �@X�Ћ��D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M���@Qh�� �M��@8�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M��E�    �E�    Q���   �M�Q�@$�СD��M�� �@Qj �M����   �СD��M�Q���   � �СD��M�Q�@�@�Ѓ����  ��� �d$ ����  �D����E�P�I�I�ыD���j ������DIj�P�E�P�A�Ѓ����5�  �D����E�P�I�I�ыD��A�M�QV�@�СD��M���@�@<�ЋD�j�j��Q�M�QP�M�BL�СD��M��P�E�P������P�B8�СD��M�Q�@�@�СD��M�Q�@�@�СD����@WS�@p�M��Ћ��h�  ��C��������]��u�E��M�j j
Q�u�@�u�p��� ������~R���� u�M����[�M��! ��_^��]� �D��M�j V�P��'  P�Bl�Ћ���jV������M�V����[�M��W! ��_^��]� �������������U���E�� �E� �E�r� �E� ]����������V���vP�N ���j ���YJ ^� �����U�������E��� �$�$��]��U���0VW��M�hTCAb�y  �M��Q  ����J �D�Phdiem�Q�M�B4�СD��M�j havem�@�@4�ЍE��E�    P�vX���E�    hsuom�KK �D��M�j hxvpi�@���   �ЉE��MСD�j hyvpi�@���   �ЉE��΍E�P�E�P�R �D��M�j haqpi�@���   �ЋD���j havpi�Q�MЋ��   �҅���   �D��M�j hrdem�@�@4�ЍE��P�I fnM���fnE���P�ǋ΃���P���W�����vX���f���7��j ����H j �h ���FX    ��j �%J �dfnM���fnE���P�ǋ΃���P���W�����vX���f���4��j ���qH �D��M�jhrdem�@�@4�ЍE��P��H �M��� �M��� _^��]� ������������ ��������VW��� �ȅ�t5�D�h-� Q�@L���   �ЋЃ���t�D�j R�A@�@8�Ѓ��3��wP����������t1j ����  ��t��趫  �؋��@P�i�  �wP���o�  ����u�j ���G _^��������������U��W�u���O�/  �u�O�$  �   _]� ����������U���HS�]���E�VW��u�����؅�u3��  贸���u�E�I% ��������  �D�S����@V�@�СD��MVQ�@�@�Ћu��E؃���P�  �D��ЋA�MQR�@�СD��M�Q�@�@�Ѓ��E��P葭  S���i�  �D�W��Mj hM  �@fE؋��   �Ѓ� ��   Ht����   E(E��   �Eȋ�P�J�  ����Y���M��H�E��Y��P�M����  �E��X �E��@�XE��E��E��E��E��E��E��E��E��E��%W�(��M���U�E�(�����E��M��oE؃��ϋ�� ��  �}  tjj j��蘬  �D��NW���   �@h�ЋM$��tIj Wj,�#� �D��M�Q�@�@�СD��M�j j�h̶�@Q�@�СD��M�Q�@�@�Ѓ��D��EP�I�I�у���_^[��]�0 ����U����} SVW��t5�K��t.�D����   �@X�Ћ���t��j ����  �����  ����u�h*� ��" ��������   �D�����IV�I�ѡD��MVQ�@�@�Ѓ��E���P��  �D��ЋA�MQR�@�СD��M�Q�@�@�Ѓ��E��P���  �} t	j�����  �D��KW���   �@h��j Wh�� � �D��MQ�@�@�Ѓ���_^[��]� ������������U��E��x;A,}�E��x;A0}	�   ]� 3�]� ������U��V�u���һ  �N<��t�f� �F<    ^]� ����������U��V�u��袻  �N4��t�D��@ �@T���F4    ^]� ��U��]�w�  �������U���SV��N��t:�D����   �@X�Ћ؉]���t!��    ���Y�  ��u#����  �؉E���u�E^[� ����3���]� ��t�WS��3��s����؅�tU�D�j S�A@�@8�Ѓ��E�3��d$ ���V�R\��tV��茤  ;Eu;}t.G�E�F��c|��u����ޣ  �؅�u��E_^[� ����3���]� �E_�0��^[��]� ����U�����W��Mf(��\}L���   f(�f(ύI �t�Y���t
f(��Y���f(ϸ   f(�t�Y���t
f(��Y����ML�   f(�t�Y���t
f(��Y����ML�   f(���I �t�Y���t
f(��Y����ML�   �Y ��Ym�YU<�M�f(��Y ��M��M��E��Y��Y��YM�YE,�X�f(��X��X��	f(ύd$ �t�Y���t
f(��Y���   f(㐨t�Y���t
f(��Y����uL�   f(�f(Өt�Y���t
f(��Y���   �t�Y���t
f(��Y����E����M��Ym�Y]D�Y��Y��YE$�YM4�X��X��X��A��]�L �������̋IV3���t"�D����   �@X�Ѕ�t����F�h�  ��u��^�U���`SVW�u���=��������D���W�@�@�СD��MWQ�@�@�Ѓ��E���P�8�  �D��ЋA�MQR�@�СD��M�Q�@�@�СD��]S�@�@�СD��MSQ�@�@�Ѓ��E   ��I ��tj���ա  �D����E�P�I�I�ыD��A�M�QW�@�СD��MЃ��@S�@x�Ѕ�tD�u����  ���MСD�Q�@�@�Ѓ���u��D��EP�I�I�у���_^[��]� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M��uQ�@�@(�ЋD����E�P�I�I�ыD��A�M�QW�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�MQ�@�@�СD��M���8�@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�СD��M��@�@Q�M�Q�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�SQ�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M��EQ�@�@�Ѓ���������U���`S��VW�K��u3���D����   �@X�Ћ�D������@W�@�СD��MWQ�@�@�Ѓ��E���P�e�  �D��ЋA�MQR�@�СD��M�Q�@�@�СD��]S�@�@�СD��MSQ�@�@�Ѓ��E   ����tg����  �D����E�P�I�I�ыD��A�M�QW�@�СD��MЃ��@S�@x�Ѕ�tA����  ���MСD�Q�@�@�Ѓ���u��D��EP�I�I�у���_^[��]� �D��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M��uQ�@�@(�ЋD����E�P�I�I�ыD��A�M�QW�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�MQ�@�@�СD��M���8�@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�Q�@�@�СD��M��@�@Q�M�Q�СD��M����@�@<�ЋD�j�j��Q�M�QP�M��BL�СD��M�SQ�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M��EQ�@�@�Ѓ������������U��V�uW�u���uV�z�  �D�V�@@�@,�ЋD������Q��jh�  ���   ��������G4�D��$h�  �A�΋��   ���_8_3�^]� �������U��V�uW�u���uV���  �D�V�@@�@,�ЋD���� �Q�$�A��h�  ���   ��� ����_8�D����$h�  �@���   ���_@�D���jh�  �@���   �ЉGH�ΡD�j h�  �@���   ��������GL�ΡD��$h�  �@���   ���_P�D���jh�  �@���   �ЉGX�ΡD�jh�  �@���   �ЉG\3�9GHt
�G8�G@_^]� ������U���0V�uW�u���uV�Ǯ  �D�V�@@�@,�ЋD������Q��jh�  ���   �҉Gh�M�D�W�QfE�M��E��@h�  Q�΋��   ��jh�  ���o �G8�~@f�GH�D��@���   ��( ��M�Gl�D�fE�Q����M��E��@h�  Q�΋��   �Ѓ����o �GP�~@f�G`�D�����$h�  �@���   ���_p_3�^��]� �������������U���0W�u���u�u虭  �D��u�@@�@,�ЋD���W���fE��E��A�M�Qh�  �MЋ��   Q�����o �G8�~@3�f�GH_��]� �����������U��V�uW�u���uV��  �D�V�@@�@,�ЋD������Q��jh�  ���   �҉G4�D�j h�  �A�΋��   ��h!D h�  �ΉG8�l �G<_^��t�u���Yy ��t3�]� �����]� ������U��V�uW�u���uV�z�  �D�V�@@�@,�ЋD������Q��j h�  ���   �҉G4�D�j h�  �A�΋��   �ЉG83�_^]� �����U��S�]VW�u���uS�	�  �D�S�@@�@,�Ѓ��E�G4    �   V����  ��t�w4F��
~�D��]��jh�  �@���   �ЉG8���D�W����$�@h�  ���   ���_@�D���jh�  �@���   ��h�e h�  �ˉGH� �GL3�_^[]� �������U��V�uW�u���uV�:�  �D�V�@@�@,�ЋD������Q��jh�  ���   �҉G4�D�jh�  �A�΋��   �ЉG8�ΡD�jh�  �@���   �ЉG<�ΡD�j h�  �@���   �ЉG@�ΡD�jh�  �@���   �ЉGD�ΡD�jh�  �@���   �ЉGH3�_^]� �����U��V�uW�u���uV�Z�  �D�V�@@�@,�Ѓ�����h�e h�  �� ������G4�D��$h�  �A�΋��   ���_8_3�^]� U��V�uW�u���uV��  �D�V�@@�@,�ЋD����X�Q�$�Q��h�  ���   ��� ����_8�D����$h�  �@���   ���_@�D���jh�  �@���   �ЉGP�ΡD�jh�  �@���   �ЉGT�ΡD�jh�  �@���   ��h�f h�  �ΉGX��
 �G\��tk���t� ��~`�O\3��f� ��~R���D��ϋ��   �@T�ЋO\VP�d� ��u#�O\V��� ��t#�D�jW�@H���   �Ѓ��O\F�� ;�|�_3�^]� ��������U��V�uW�u���uV芨  �D�V�@@�@,�ЋD�����Q�$�Q��h�  ���   ���_8�D���W��΋@�$h�  ���   ���_@�D���j h�  �@���   ��������GH�ΡD��$h�  �@���   ���_P�D���jh�  �@���   �ЉGX3�_^]� ��U��S�]VW�u���uS詧  �D�S�@@�@,�ЋD������Q�$�Q��h�  ���   ���_8�D���jh�  �@���   ��h�f h�  �ΉG@�� �GD��tl��蕕 ��~a�OD3�臕 ��~S�I �D��ˋ��   �@T�ЋODVP脔 ��u#�ODV�� ��t#�D�jW�@H���   �Ѓ��ODF�4� ;�|�_^3�[]� �������U��V�uW�u���uV誦  �D�V�@@�@,�ЋD�W�Q���$h�  �Q�΋��   ���_8�D���W��΋@�$h�  ���   ��������_@�D����$h�  �@���   ��������_H�D����$h�  �@���   ��������_P�D����$h�  �@���   ��������_X�D����$h�  �@���   ���_`_3�^]� �U��V�uW�u���uV芥  �D�V�@@�@,�ЋD�����Q�$�Q��h�  ���   ���_8�D���j h�  �@���   �ЉG@3�_^]� �������������U��V�uW�u���uV�
�  �D�V�@@�@,�ЋD������Q�$�Q��h�  ���   �������_8�D����$h�  �@���   ���_@�D���W��΋@�$h�  ���   ���_H�D���jh�  �@���   �ЉGP3�_^]� ��������������U��V�uW�u���uV�:�  �D�V�@@�@,�ЋD�W�Q���$h�  �Q�΋��   ���_8�D���W��΋@�$h�  ���   ���_@�D���W��΋@�$h�  ���   ���_H�D���j h�  �@���   �ЉGP���D�W����$�@h�  ���   ���_X�D���W��΋@�$h�  ���   ���_`�D���W��΋@�$h�  ���   ��������_h�D����$h�  �@���   ���_p�D���j h�  �@���   ��������Gx�ΡD��$h�  �@���   ��ݟ�   _3�^]� ������U��V�uW�u���uV蚢  �D�V�@@�@,�ЋD���� �Q�$�Q��h�  ���   ���_8�D���jh�  �@���   �ЉG@3�_^]� �������������U��V�uW�u���uV��  �D�V�@@�@,�ЋD������Q��j h�  ���   �҉G4�D�jh�  �A�΋��   �ЉG8�ΡD�j h�  �@���   �ЉG<���D�W����$�@h�  ���   ��������_@�D����$h�  �@���   ���_H�D���W��΋@�$h�  ���   ��������_P�D����$h�  �@���   ���_X�D��@��������   ���$h�  ���_`�D���W��΋@�$h�  ���   ��������_h�D����$h�  �@���   ��������_p�D����$h�  �@���   ��������_x�D����$h�  �@���   �������ݟ�   �D����$h�  �@���   ��ݟ�   _3�^]� ��������������U��V�uW�u���uV��  �D�V�@@�@,�ЋD�����Q�$�Q��h�  ���   ���_8�D���W��΋@�$h�  ���   ��躾 �G@�ΡD�jh�  �@���   �ЉGD3�_^]� ���U��V�uW�u���uV�J�  �D�V�@@�@,�ЋD������Q��j h�  ���   �҉G4�D�j h�  �A�΋��   �ЉG8���D�W����$�@h�  ���   ��������_@�D����$h�  �@���   ���_H�D���jh�  �@���   �ЉGP3�_^]� ����������U��]�w�  �������U��V�uW�u���uV�Z�  �D�V�@@�@,�ЋD������Q��j h�  ���   ��������G4�D��$h�  �A�΋��   ���_8_3�^]� �������U��SV�uW�u���uV�ٝ  �D�V�@@�@,�ЋD�����Q�$�Q��h�  ���   ���_8�D���W��ˋ@�$h�  ���   ���_@�D���jh�  �@���   �ЉGH3���L�D���j �P��M  P���   ��F����|�_^3�[]� �����������U��V�uW�u���uV�
�  �D�V�@@�@,�ЋD�����Q�$�Q��h�  ���   ��������_8�D����$h�  �@���   ���_@�D���j h�  �@���   �ЉGH3�_^]� ���U���u�u�u�o�  3�]� ���������U���0V�uW�u���uV�G�  �D�V�@@�@,�ЋD������Q��j h�  ���   �҉G4�D�jh�  �A�΋��   �ЉG8�ΡD�j h�  �@���   �ЉG<���D�W����$�@h�  ���   ���_@�D���W��΋@�$h�  ���   ��������_H�D����$h�  �@���   ��������_P�D����$h�  �@���   ��W��_XfE�D��M�Q�E��M�h�  �@Q�΋��   �ЍM�Qh�  �o �M�Q�G`���~@f�Gp(0��D�fE��p��E��@���   �ЍM�Qh�  �o �M�Q�Gx���~@fև�   W��D�fE��E��@���   ��jh�  ���o ���   �~@fև�   �D��@���   �Љ��   3�_^��]� �����U��V�uW�u���uV�*�  �D�V�@@�@,�ЋD������Q��j h�  ���   �҉G4���D�W��$�A��h�  ���   ��������_8�D����$h�  �@���   ���_@�D���jh�  �@���   �ЉGH�ΡD�jh�  �@���   ��h�e h�  �ΉGL��  �GP3�_^]� ������U��V�uW�u���uV�:�  �D�V�@@�@,�ЋD������Q�$�Q��h�  ���   ���_8�D���jh�  �@���   �ЉG@�ΡD�jh�  �@���   �ЉGD�ΡD�jh�  �@���   ��h�f h�  �ΉGH�L�  �GL��tu���� ��~j�OL3���� ��~\�
��$    �I �D��ϋ��   �@T�ЋOLVP�ԅ ��u#�OLV�g� ��t#�D�jW�@H���   �Ѓ��OLF脆 ;�|�_3�^]� ��������U��V�uW�u���uV���  �D�V�@@�@,�ЋD������Q��j h�  ���   �҉G4�D�jh�  �A�΋��   �ЉG8�ΡD�jh�  �@���   �ЉG<3�_^]� ���������U��V�uW�u���uV�j�  �D�V�@@�@,�ЋD����X�Q�$�Q��h�  ���   ��� ����_8�D����$h�  �@���   ���_@�D���W��΋@�$h�  ���   ���_H�D���jh�  �@���   �ЉGP�ΡD�jh�  �@���   �ЉGT�ΡD�jh�  �@���   ��h�f h�  �ΉGX�-�  �G\��ti���τ ��~^�O\3���� ��~P�D��ϋ��   �@T�ЋO\VP��� ��u#�O\V�T� ��t#�D�jW�@H���   �Ѓ��O\F�q� ;�|�_3�^]� �����U��W�u���u�u��  �D��u�@@�@,�ЋD����ЋA��j h�  ���   �ЉG43�_]� ���U��SVW�u�}���uW處  �D�W�@@�@,�ЋD����ϋ����   �RT�ҋD�hK  Ph�  �Q�΋Bl��h.� P�C4�q������t_^�����[]� �K4��t�D��u�@ �@P��_^[]� _^3�[]� U��V�uW�u���uV���  �D�V�@@�@,�ЋD������Q��j h�  ���   ��j h�  ��fn�����G8�D��@���   �Ѓ���fn�����G@W��D��$h�  �@���   ���_H�D���W��΋@�$h�  ���   ���_P�D���W��΋@�$h�  ���   ��������_X�D����$h�  �@���   ��������_`�D��$h�  �@���   ����������_h�D����$h�  �@���   ��������_p�D����$h�  �@���   ���_x_3�^]� �����������U��} SW�}��tM�K��t6�D�V���   �@X�Ћ���t��3���;���P�!�  ���j�  ����u�^j Wh�� �� ���D��KW���   �@h��_[]� ��������̋A�������������U����}u{V�u��    tm�E��E�  P�E��E�    P�E��P�E�P�E�P��U ��u�����ȉE��M��M��E��M��P�E�P�H �M�E�j j�j QP���   �����^��]������U��}uj h�� �;� ��]�������U����}u|V�u�E�P�E��E�  P�E�E�    P�E���P�E�P�'U ��u�����ȉE�Q�M���   P�)���^��]ËM��E��M��P�E�P��G �M�E�QP���   �����^��]�����U���  VW��� t�u�u�u�uV��  ��_^��]� �u��j �u}  j�ΉE�i}  j�ΉE��]}  �MW��E�W�f(�����m����E�fM�fM�fM�fM���tL�D�j Q�@@�@8�Ѓ���l�����u�u�uQ�ȋBH���m�W��o fE�fE��~@�E��M���tD�D�j Q�@@�@8�Ѓ���l�����u�u�u�Q�ȋBH���o�~hfM�fM��m�� ��   ����   �D�j V�@@�@8�Ѓ���l�����u�uVQ���RH�GH��wu�$�����l����4��t����*��|���� ��t����X�l����X�|����Y��W��M�f/�v
(��M�����f/�v(��M���M����� �m�t�\�(��M�fMЋG4W�HfEȃ���  �$���fE��]��E�f��  �E�f/�vf(��f(��M��u�f/�w(��E��}�f/�w(�f��E��A  �}�f(��u�f(��YM�(��YE��Ye�f��M��  fE����]��ă��f�h��� f�X��l���P��Q���o ��4�~`�E��  fE����]��ă��f�h��� f�X�E�P�qR���fE����]��ă��f�h��� f�X�E�P�R����E�f/�vf(��f(��U��M�f/�w(��E��}�f/�w(�f��E��  fE����]��ă��f�h��� f�X������P�SS������fE����]��ă��f�h��� f�X��$���P��S��������}�f(��u�f(��XM��Xe�(��XE�f��M��|  fE����]��ă��f�h��� f�X��4���P�ST���h���fE����]��ă��f�h��� f�X��T���P��T���1���fE����]��ă��f�h��� f�X��d���P�UV�������fE����]��ă�� f�X���f�h������P�~T�������fE����]��ă��f�h��� f�X�����P�WX������fE����]��ă��f�h��� f�X������P��Y���U���fE����]��ă��f�h��� f�X��<���P��Z������fE����]��ă��f�h��� f�X�����P�\��������U��}��M��\��u��P��\��e��\�fT�fT�f�fT��U��}  �E�f(��]����X��u��Y�(��}��YE��\��E��X��Y��Y��\��E��X��Y�f��Y��]��\��  �}�f(��u�f(��\M��\e�(��\E�f��M���  fE����]��ă��f�h��� f�X������P��]�������fE����]��ă��f�h��� f�X������P�?^������fE����]��ă��f�h��� f�X��|���P�^���]���fE����]��ă��f�h��� f�X��L���P�Q_���&���fE����]��ă��f�h��� f�X�����P�^�������fE����]��ă��f�h��� f�X������P�c_�������}�f(��u�f(��\U����f(��\M��\e��X��X��X�f��U��Q�}�f(��u�f(��XU����f(��XM��Xe��\��\��\�f��U��W��}��u��U��M��\��]��\��E��\�E�Y��Y��Y��G8�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� ��������e�}�����@�q�����"�Y�������0�g������C�����(�_������;�r���������������U������$  SVW��� t�u�u�u�uV�G�  ��_^[��]� �Mj �s  �M��j�\$�s  ������L$��u�EW� �@_^[��]� � �]��   ����   �D�j V�@@�@8�Ѓ��L$x��uSVQ���RH�GH��wx�$����T$x�6��$�   �+��$�   � ��$�   �XT$x�X�$�   �Y�����W�f/��T$v(��T$�"f/�v(��T$��T$W����� tf(��\�f(��T$�WۋGL�   �\$0W��\$8�щL$�T$f�$�   ;�wU�$����L$�T$�D�   �щL$�T$�3�   �щL$�T$�"�OX���L$%  �yH���@uA�L$�щL$�O8fn�����D��t$j V�@@�^ȋ@8fn�����L$x�O@�^��L$h�Ѓ��L$H��uSVQ���RH�O8W�f.��o �~X��\$h�d$x��$  ��Dz*�\ �   �t$�T$pt�E� f�X_^[��]� �t$�G@f.��Dz�D$   �T$`f.ʟ��Dz
f.��D{���$�   W�f�$�   f�$�   f�$�   f�$�   ��tjh��$�   SP��� ���L$����  ��$�   �A���$�   ��$�   ��$�   �\$`�+��d$ �����l$(�D$@fn�����Y��X���$�   ���  �L$�F��+L$D�������	��$    ����$�   �\Cfn�����Y��YT$p�X���$�   �\K��$�   �\�Y��Y��X��X�輽 �G\f(ȃ� ��   H��   H�Q  �G8f/��B  �^ȡD�j �@@�@8����t$�\���$�   �Ѓ���$�   ��uQ�t$�L$TQ���RH��$�   �D$H�L$P�T$X�Y��Y��Y��XD$(�XL$ �X\$8�XT$0f(�f(��l$(�d$ �T$0�\$8�   �G8f/���   �D�j �t$�@@�@8�Ѓ���$�   ��uQ�t$�L$TQ���RH�D$H�XD$(f(��D$P�XD$ �l$(f(��D$X�XD$0�d$ �D$0�D$8�X���D$8��d$ �l$(�F�L$D�"����\$`�t$�L$�D$@�S@I�D$@�L$������D$8W�f/�v(����^��t$h(�(��YL$0�Y��Y��+�oD$x�t$h��$�   ��$�   f���$�   �  ��$  u(Ճ$ ��$   u(܃( u(��D$�\��\܋E�\��Y��Y��Y��GP�X��X�_�X�^�\��\�[�\��Y��Y��Y��X��X��X�f��f�H��]� ����������������U���PVW��� t�u�u�u�uV莂  _��^��]� �MSj ��l  �M��j��l  W�W��E�������E�fM�fM���t=�D�j S�@@�@8�Ѓ��Mȋ�u�uSQ���RH�o fE�fE��~@�E�� [��   ����   �D�j V�@@�@8�Ѓ��Mȋ�u�uVQ���RH�GH��wc�$�\��E��%�E���E���E��XE��XE��Y��W��E�f/�v
(��E�����f/�v(��E���E����� t�\�(��E��h fE��m��u�f��E�tE�  t�_8f/�w�]ȃ$ �U�t�G@f/�v(Ѓ( t�GHf/�v(��
�U��]ȃl t<�  t�GPf/�v(؃$ t�GXf/�v(Ѓ( t�G`f/�v(��M��\��E��\��\�E�Y��Y��Y��Gp�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� �I ������������U��y t�u�u�u�u��  �E]� �oA8�E� �~AHf�@]� �����U���hVW��� t�u�u�u�uV�  _��^��]� �Mj �
j  ��W�WɅ��^  �D�j V�A@�@8�Ѓ��M���u�uVQ�ȋBH�ЋO4����~H�o �E�����   �$�h��o �E��~@�E�P�E�f�E�P�>� �Mȃ��{�o �E��~@�E�P�E�f�E�P�� �M����Q�o �E��~@�E�P�E�f�E�P�� �M����'�M�� �M���E��XE��X��Y��(ȋG8�M�Ht3HuB�E����� ����]��E��\�fTP��\���E���軛 �]��M��O<�E����$P�I �o �~H�E_^� f�H��]� B�l���������U���xVW��� t�u�u�u�uV��}  ��_^��]� �Mj �:h  ��W��E�W�fE���]  �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�O4���ofE��~J�M�;O8�  It_It(Iu|�o����� �~Bf�@�E�P�qT�����D�o�E�P�EЍE��~BPf�E��� �oE����~M�fE���E�P�E�P�ۖ ���o fE��~H�M��G8HtZHtHur����� f�H�E�P�rU�����H�E�f�M�P�E�P�E��Ɨ �E���oE��~M�� f�H_^��]� �E�P�E�P�H� ���o fE��~H�E� f�H_^��]� �E_^�f�@��]� ���������������U���   VW��� t�u�u�u�uV�|  _��^��]� �4 W�W�u�E_^�f�@��]� S�]��j �Df  �����  �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�G8�������   �$�p��oE��E�P�EЍE��~E�Pf�E�莖 �E����   �oE��E�P�EЍ�p����~E�Pf�E��]� ��x������W�oE��E�P�EЍE��~E�Pf�E��/� �E����,�E��%�E���E���E��XE��XE��Y���OL�E����$P�N ���W��Hf/�v(��	f/�v(ʋw4f(�f.�fn������^���Dz����   �E��   f.ʟ��Dz(��   3���~2��I fnЍH���fn�����Y��Y�f/�rf/�w��;�|�W�E[_^� f�X��]� ���p�L$�D$�$��3�������%���]��E��E���~��G@��f.�V���DzN�,d  ����u�EW�[_^� f�@��]� V�x}���M���Q�MQV�M�Q���RH�o �~X�S���W��]�fE�f(��E�W�fE���c  �E��t4P�#}���M���Q�MQ�u�M�Q���RH�o �~Xfe��]���]�W��M�W�f/���   �o@�\�f.���D{�X���\��^�(����$�X0�����]���u�H t�w4��e�f�]��AN��~<V���	c  ����t.V�m|�����M���u�uVQ���RH�o �E��~@�E��U��Y���M��\M��]��X���\]��Y��Y��XM��X]�f(��M��\M��Y��XM�f���������f(��\o@�\�f.П��Dz(���\��^ʃ��$�a/���G4���]�;�u�H tj��e�f�]��AF;�<V���b  ����t.V�u{�����M���u�uVQ���RH�o �E��~@�E��U�W��Y���M��\M��]��\]��X��Y��Y��XM��X]�f(��M��\M��Y��XM�f�������I ���P�{�������������U���0VW��� t�u�u�u�uV��v  _��^��]� �Mj�*a  ����u�EW�_^ �@��]� �D�j V�@@�@8�Ѓ��M��u�uVQ���RH�Mj ��`  ����u�E�oE�_^� �~E�f�@��]� �D�j V�@@�@8�Ѓ��MЋ�u�uVQ���RH�4 �M��U��E�t!�G@�� tHt
Hu�M���U���E�8 t!�GD�� tHt
Hu�M���U���E��< t�GH�� t)Ht!Ht�M��E�oE�_^� f�H��]� (���(����������������U���pVW��� t�u�u�u�uV�^u  _��^��]� �MSj �_  �M��j�_  ���W��M����E�fM�fM���t=�D�j S�@@�@8�Ѓ��M���u�uSQ���RH�o fE�fE��~@�E�� [��   ����   �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$����E��%�E���E���E��XE��XE��Y��W��E�f/�v
(��E�����f/�v(��E���E����� t�\�(��E��  fE��E�t �E��E��O4���$P�G �@��E؃$ �E�t �E��E؋O4���$P�G �@��E��( �E�t �E��E��O4���$P�_G �`��~e��oUȋE�u��m��\��]��M��\��E��\��Y��Y��Y��G8�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� �������U���(  VW���}�� t�u�u�u�uV��r  ��_^��]� �uW�W��~T ��  �Mj �]  ( �������U��M�f�8�����tA�D�j R�A@�@8�Ѓ���������uV�u�Q�ȋBH���o ��8����~@�E��P W��NTfE��E��o��   �E��~��   f�E��o��   �������~��   fօ ����o��   ��P����~��   fօ`���u�o��   �E��~��   f�E�3�9��  Q��3�9WTD�3��E�D��}��@�@X���Mȃ��E����J  �M��E�D�W�vT�@�@T�Ћ����E��x\ t>�D����   �M�RT���wP�E��H\��[ �M�3�9QX��3Ƀ����;���  �vTW�j �D�j�o��   ��@  ������~��   fօ���W�f�p����M�fE��M���(  ���   Q�u��@��P�����RQ��d  ������Q�M�Q�����Q�M�Q��p���QWV�Ћu��8���  ���  �E    �E�    �9 t$�E�P�EP�FT��0  Q誒 ���} ��  ���   W�W�f(�u}�D�W��VTfE��M�f� �����0����H�� ���P�E�P��(  ��P���P�E�P�����P���   ��P��`  ���$jj WR���oe���4�~]��   �E��YE��FT�U��YU��X��E��YE��X���  �Y�f/�rZ��8  f.����D{4fTP�fW`���h����c� f(���h����"� f(��f(�fTP�f(�f�}��� ���G@�D$� f�X�� ���P�+���G8��$�o�~X�Y]�f������������Y�p����Y�x����Y��Y��Y�W�f/�v(�f/�v(�f/�vf(��E��X��E��E��X��E��E��X��EءD��}��vTG�@�}��@X�Ѓ�;�������E��M��Y�8����Y�@���f(��E��YE�fыE_^�f�@��]� ���U����   VW��� t�u�u�u�uV��m  _��^��]� �u��j �%X  j�ΉE�X  ������M�E���u�EW�_^ �@��]� � ��   ����   �D�j V�@@�@8�Ѓ��M܋�u�uVQ���RH�GH��wd�$����M��%�M���M���M��XM��XM��Y��W��M�f/�v
(��M��f/��v����M���M�� �Mt����\�(��M��GH�   W�W��U�fE�;�w)�$����   ��   ��wX��%  �yH���@uF�O8fn�f(����f.��^؟�]���Dz
�   �U��D�j Q�@@�@8�Ѓ��M���u�u�uQ�ȋBH���o ��|����~@�E�E�W���T���f����f�$���f�4���f�D�����tjhP�����P�T� ��3��E���)  �E��E��E��E��G@fW`�fn�����E��YM��M��� �YEċE�X ������E��ɑ �YEċEj �u�X@�D�������@@�@8�Ѓ��������uQ�u�M�Q���RH�E��XE�E�@�E�f(��E��XE��U�f(��E��]��XE�f(��e�;��/�����~Ofn�W����f.���D{����^�(��Y��Y��Y��f(�f(�f(���]��U��eԃ  ��|���uf(Ճ$ �M�uf(ك( �u�uf(��E��\��\ًE�\��Y��Y��Y��GP�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�`��]� ��J�Q�X�_��������U������  ��3ĉ�$�  �ES�]V�uW���D$D� t�uSPV�i  �  �CTW�WɅ��g  fD$x�D$p    f�$�   �D$l    f�$�   Ǆ$�       f�$  f�$   f�$0  f�$@  f�$P  f�$`  f�$p  f�$�  f�$�  f�$�  ����$�   ��$�  ��$  ���   �T$0���   ���   (��Y��L$H(��Y��\$8�X�(��Y��X�負 f(�W�f.џ��DzW��L$`fD$P�<����^��L$0�T$8�\$H�Y��Y��Y��L$X�T$`�\$P�D$PP�CT���   ��P��$�   P�x �KT�T$t������D���$  �o��   R�T$4��$�   R�~��   ��$�   ��$H  ���D$D    ��$8  �D$@    ��$   �o�$�   fք$�   fք$`  fք$H  fք$0  �~�$�   fք$  fք$�  fք$�  fք$x  �G8��$   ��$�  ��$�  ��$h  �@�$RQ��$  �Ѓ���uW��f�F��   �|$4�t�D tP�D$h�D$8��tD���    t;�D��L$D���   �@T�ЋL$8���   �ODP�[Q 3�9W@��3Ƀ����;�t��CT���   ���   �\�$�   �\T$x���   �\�$�   �Y��Y��Y��X��X��k� �^G8���W��\�f/�w(�f(�f��f�N��$�  ��_^[3��:� ��]� ����U����   VW��� t�u�u�u�uV�e  _��^��]� �u��Sj �P  j�΋��	P  j�ΉE��O  ����E��E����  �D�j S�A@�@8�Ћu�M�����uVSQ���RH�M�~H�M��o �E�����  �D�j Q�@@�@8�Ѓ��MЋ�uV�uQ���RH� �o �E��~@f�E���   �E����   P�h���M����uVQ�M�Q���RH�GH��wc�$�<�E��%�E���E���E��XE��XE��Y��W��E�f/�v
(��E�����f/�v(��E���E����� t�\�(��E��WHW��_PW���X����^8��^8��U��]�f����f�(���f�8���f�H�����tjh�����VP�g� �U����]�W��%��f.џ��Dz
������'�E��\��^��YGX�X�����\G8�����f.ٟ��Dz
�� ����'�E��\��^��YGX�X� ����XG@�� ����D�j S�@@�@8�Ѓ��������uQS�M�Q���RH�  �u�uf(���M��$ �e�uf(���]��( �m�uf(���U��E��\��\܋E�\�[�Y��Y��Y��G`�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�P��]� �E[_^� f�H��]� �EW�[_^ �@��]� �I ������������U������L  �y SVW�L$@t�u�u�u�uV�b  ��_^[��]� �Mj �`L  W�Wɋ��L$ �L$p�L$0fD$`fD$HfD$`��u�E�H_^[��]� �M��$�   f�$�   f�$�   f�$�   ��tjhQ��$�   P�� �M���D$P����\$`�D$(�D$H�D$H�D$h�T$D�D$8�\$�d$ �D$@�4�    fn������Y@8�XA��$�   ��$    fn�����Y@8�@@�X�D$x�� ��  H�  H�  9�X���   �D�j S�@@�@8��fn�X���$�   �������u�D$QS�L$lQ���RH�\$�H�P� �Y��Y��Y��XL$(�XT$ �\$�XD$H�L$((��L$ �D$H��|� �p  �D�j S�@@�@8��fn�|���$�   �������u�D$QS��$4  Q���RH�\$f(��Y �H�P�Y��XD$�Y�f(���  ��� ��   �D�j S�@@�@8��fn����$�   �������u�D$QS��$L  Q���RH�\$� �H�P�Y��Y��Y��XD$H�XL$(�\$�XT$ �D$H�L$(�T$ ��4� �]  �D�j S�@@�@8��fn�4���$�   ���uQ��$�   ��   ���� ��   �D�j S�@@�@8��fn�����$�   �������u�D$QS��$  Q���RH�\$f(��H�P�Y �Y��Y��XD$H�XL$(�\$�XT$ �D$H�L$(�T$ ��� ��   �D�j S�@@�@8��fn����$�   ���uQ��$  ����SQ���D$ �RH�\$� �H�P�Y��Y��Y��XD$(��XL$8�XT$0�\$�L$8�T$0�D$@G�M����������T$DB�T$D���f����D$H�Y��Y��X�迕 �L$(�D$H�D$8�Y��Y��X�蜕 �L$0�D$�D$ �Y��Y��X�(��v� fT$H�E�L$_f�^�[f�@��]� �U����   VW��� t�u�u�u�uV��\  _��^��]� �MSj �FG  �M��j�:G  ������E�����  �D�j S�A@�@8�Ѓ��M���u�uSQ���RH�o �E��E��~@�E�E�W���h���f�(���f�8���f�H���f�X�����tjhP��(���P�ė ���GH藒 �YG@�X�(�����(����GH�x� �YG@�D�j S�X�0�����0����@@�@8�Ѓ���(�����uQS�M�Q���RH� �o �E��~@�E���   ����   �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$��	�E��%�E���E���E��XE��XE��Y�����W�f/��E�v
(��E�� f/�v(��E�����W��E�� t�\�(��E��W�  �oE��}��u�f��E�t$�P tf(��f(��M��\��YO8�X���M��$ �m�t$�P tf(��f(��U��\��YW8�X���U�( t�P t(��]��\��Y_8�X��E��\΋E�\��\�[_�Y�^�Y��Y��X��X��X�f��f�X��]� �EW�[_^ �@��]� %��������U���   VW��� t�u�u�u�uV�Y  ��_^��]� �u��j �D  j�ΉE�	D  ������M�E�W����  �D�j Q�@@�@8�Ѓ��M���u�u�uQ�ȋBH�Ѓ �o �~H�E��E��M���   ����   �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$���M��%�M���M���M��XM��XM��Y��W��M�f/�v
(��M�����f/�v(��M���M����� t�\�(��M��oE��E�P�EȍE��E�Pf�E��(q �G8���P �^@�t�E��G@�E��M�XE��E��E����u �E�W��O@�Y���Y��]��X���\��Y��X��M��E�P�E�P�q �wHW��f/��o �E��~xv�%��f(�f(�f(��fT5P�f(�f(�f(��%���\U��\]��\���ă��Y��Y��Y��XU��X]��X�f��WX(�(��]��XE��XM��X�f�����f�P�E��D$�G`�X��U��M��$P�x�������o �E��~@f�E����   �D$�o ��~@�E�Pf�A�����$�x �o �E��~h�]�tR�OhW�f/�v(��e�f/�v(�f/�v(��Opf/����v(�f/�v(�f/�v
(���e��\]��\e��\m��U��E�Y��Y��Y��X]��Xe��Xm�f��f�h_^��]� �EW�_^� f�P��]� ���
�
�
�
����U������@�y t�u�u�u�u�U  �E��]� �U�BT��u����\B���^  �y@ �o��   �~��   �D$(u�o��   �~��   �D$(���   W��-`��T$0�|$(�@ �XfW��H(fW��Y�fW�f(��Y��X�f(��Y��X�f/����v
����f(��L$0�X �Y�fW��Y��Y��A8�L$�H�Y\$fW��Y��Y��$�@(fW��X��Y�f(��-���X�f(��\$ �Y��P��\��$�\�(�fT�f(��\��X��Y��Y�f.��L$�T$���Dz�d$�#(�fT��Z� �L$W��P��D$f.̟��Dzf(��fT�f(��&� f(�W��\$ f(��X��Y��XL$f.̟��D{1�|$f(��Y,$f(��Y�f(��X��Y��X�f.ԟ��Dz!�E( �����f�@��]� �\�f(�fW`��\��Y��Y��Y��X\$�X��^��^��X��Y��f(ȋEf��f�@��]� ���U���xSVW��� t�u�u�u�uV��R  ��_^[��]� �Mj �H=  �M��j�<=  W�W��M���fE�����E���t8�D�j S�@@�@8�Ѓ��M���u�uSQ���RH�o �E��~@�E�� ��   ����   �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��w`�$�t�E��%�E���E���E��XE��XE��Y�����W�f/��E�v�M��f/�v(��M������M�� tf(��\�f(��M��W@W��OH�\�f.ȟ��Dzf(���]��\��^�f.ȟ��Dzf(���e��\��^�f.ȟ��Dzf(���u��\��^��GP�� �WX���\�f(�(��Y��gh�Y��Y��X��_`�X��X����Y�f�(��E�f(��Y��YE�(��X��X��X��Gp�D$f��f�`�E�P����_x��$���w4�o���o)���~a�m�� f�f�@��%���M����]��E���\���\��\��Y��Y��Y��X��X��X��P�f��(f�`�E��D$���   �$P����mЃ�,�  �o �~X�E�uf(���M��$ �u�uf(���U��( �e�u(܃8 t W�f/�vf(�f/�vf(�f/�v(؃< t%���f/�vf(�f/�vf(�f/�v(��E��\��\֋E�\��Y��Y��Y����   �X��X�_�X�^�\��\�[�\��Y��Y��Y��X��X��X�f��f�X��]� ��V]dk������������U������$  SVW���|$D� t�u�u�u�uV��N  ��_^[��]� �Mj �9  ��W��L$��u�E� f�@_^[��]� �G@�   �D$0�D$(�\$fD$h;�w1�$���   ��   ��_D�É\$%  �yH���@uC�\$�O8fn�����D�j Q�@@�^ȋ@8�L$h�Ћu��$�   ����uV�t$Q���RH�G8W�f.��o�~P��T$X��$�   ��$�   ��Dz�E�f�P_^[��]� �����$  �^�W���$�   f�$�   f�$�   f�$�   f�$�   ��tjh��$�   VP�� �����  �D$p�C���$�   ��$�   �+��D$H�D$h���ȉ\$���D$8���L$T�D$��I �\$`��fn�����Y��X��D$ ��$�   ���$    �\Ffn�����Y��Y��X���$�   �\N��$�   �\�Y��Y��X��X��Ǆ �D$D�H8f/���   �Y�$�   �D����j �t$�@@�\ȋ@8�L$(�Ѓ���$�   ��uQ�t$��$�   Q���RH�\$ ��$�   ��$�   ��$�   �Y��Y��Y��XD$8�XL$H�X\$(�XT$0f(���$�   f(��d$8f(��l$Hf(��|$(�t$0�D$ ��D$ �d$8�l$H�t$0�|$(�G�\$`K������D$�V@�L$�\$�L$T�D$�W���W�f/�v ����^��\$X�Y��Y��Y��%�o�$�   �\$X�D$h�l$pf��d$h��$�   �\���$�   �\�����\͋E_�X��X��X�^[f��f�X��]� ��C$+������������U���   VW��� t�u�u�u�uV�{J  _��^��]� �uW�f]�W��FT����   �G4���2  �$�|�=���\~�  ����g �]��F���g �]��F���zg �Ef]�_�]��}��^f�x��]� �E( ��=��_�^f�x��]� �P �o��   �~��   �E��e�u�o��   �~��   �E��e��O4���l  �$�����   �E��=���H �YM��Y@�X��@(�Y��X�fTP��\��  ��0  ���  �o��  _�~�   �E^�f�x��]� �o�  _�~�   �E^�f�x��]� �8 t&��   ���D$G@$�������  ��   �  ��0  ����  �o��   �]��o�(  ��h����o�  �U��o�8  f��Y��o�  �X��E��om�f(���0  �Y��Y��X�(�f��YE��X�f(���   �Y��m���P  �X��X��E��o�H  �8 �YE��M��Ym��Y��X��Y��X��M��oM��U����X�f��X���  ����Y��Y��Y��X��X��X�f(ًEf�_^�f�x��]� ���in���]�W��U��o@`�o��   ��h����o@p�o��   f��Y��o��   �X��E��om�f(����   �Y��Y��X�(�f��YE��X�f(����   �Y��m����   �X��X��E��o��   ������8 �o�f���   ���(��E��U��Y��Y��Y��X��X��X�f(���������   �@�H �YE��YM��X��@(�Y�3��X�f/�����fn�����$�������]��}�(�fߋE_^�f�x��]� ��;M;MMM��w���E����U���@VW��� t�u�u�u�uV�E  _��^��]� �MSj ��/  �M��j��/  W�W��M���fE�����E���t8�D�j S�@@�@8�Ѓ��M؋�u�uSQ���RH�o �E��~@�E�� [��   ����   �D�j V�@@�@8�Ѓ��M؋�u�uVQ���RH�GH��wd�$���M��%�M���M���M��XM��XM��Y��W��M�f/�v
(��M��f/��v����M���M�� t����\�(��M��-���M�f(��E��\��u�f(��e��\ЋE�\�_�\�^�\��\��Y��Y��Y��X��X��X�f��f�h��]� ������U��y t�u�u�u�u��C  �E]� �EW� �@]� �������������U���xVW��� t�u�u�u�uV�~C  _��^��]� �u��Sj ��-  j�ΉE��-  j�΋���-  �MW��E�f(��e�Wɋ�fE�����E�fM�fM���tB�D�j Q�@@�@8�Ѓ��M���u�u�uQ���RH�e�W��o �E��~@�E���t=�D�j S�@@�@8�Ѓ��M���u�uSQ���RH�o�~`fM�fM��e� [��   ����   �D�j V�@@�@8�Ѓ��M���u�uVQ���RH�GH��wc�$�`$�E��%�E���E���E��XE��XE��Y��W��E�f/�v
(��E�����f/�v(��E���E����� �e�t�\�(��E�fM؋G4f��u��m��MЃ��  �$�p$�  t�M��X���MЃ$ t�U��X���U؃( ��  �}�(��X���  �  tf(��\M���MЃ$ tf(��\U���U؃( ��  f(��\]��  �  t�M��Y���MЃ$ t�U��Y���U؃( �V  �}�(��Y��E  �  W�t)f.���D{�U�f.П��D{
f(��^��f(���MЃ$ t)f.���D{�}�f.����D{
f(��^��f(���U؃( ��   f.����D{�}�f.����D{f(��^��   (��   �  t�M�f/�v
(���MЃ$ t�U�f/�v
(���U؃( tf�E�f/��E�  t�M�f/�v
(���MЃ$ t�U�f/�v
(���U؃( t�E�f/��f���f(��
�U��M��E��\��\֋E�\��Y��Y��Y��G8�X��X�_�X�^�\��\��\��Y��Y��Y��X��X��X�f��f�X��]� 4!;!B!I!�!&"j"�"T#�#��������U����   S��V�]��{ t�u�u�u�uV��>  ��^[��]� �u��Wj �!)  j�ΉE�)  �} ������E�W�u�E_^[� f�@��]� �{ ��   ����   �D�j W�@@�@8�Ћu�Mă���uVWQ���RH�CH��wd�$��(�M��%�M���M���M��XM��XM��Y��W��M�f/�v
(��M��f/��v����M���M��{ t����\�(��M���u�D�W��}j W�@@fE��E�    �E�@8�Ѓ��������uVWQ���RH�K8�YX��M�o �M��E��~@�E�W���h���f�(���f�8���f�H���f�X�����tjhQ��(���P�x �M����U̍{L�m�3��]�U��m����    �? �  ����̋��������+�fn�����\��Y��X�(�����(���fn�����^8��E��E��$��v �]��,E�j Sfn��D�����\��YE��X�0�����0����@@�@8�Ѓ���(�����uQS�M�Q���RH�M��M��U��o�]��u���(����~A�M�fօ8����fn�����M��Y��Y��Y��XM��XU��X�(��m��U��]���]�M��M�F����������]��{H tJ��tFfn�W����f.����D{$����^�(��Y��Y��Y�f(�(��f(�(�f(���u��m��e܃{  �K@f(�(��X��m��X��X�uf(Ճ{$ �e�u(܃{( �u�u(��E��\ՋE�\��\�_^�Y�[�Y��Y��X��X��X�f��f�H��]� P%W%^%e%��������U��y Vt�u�u�u�uV�:  ��^]� �Mj ��$  ����t-�D�j V�I@�I8�у��ȋ�u�uV�uV�RH��^]� �EW�^ �@]� �������������U������(  VW���|$$� t�u�u�u�uV��9  ��_^��]� �Mj �P$  �O@���Y��W��L$�D$�D$�X ��L$0��u�E �@_^��]� �D�j Q�@@�@8��W����E���D$xfD$8fD$HfD$XfD$h��tjhP�D$@P��t ���M����\$@�T$8�t$,��    �T$$���fn�����D$(���YB8�X��D$@fn��BH����YB8�X��D$8�� ��  H��   H�R  9�X�ta�Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn�X��M����Y��XD$(��L$��|� ��  �Q�L$<Q�t$�@H��$  Q�����o�~P(�f�f/�vf(�f/�vf(�fn�|��   ��� t^�Q�L$<Q�t$�@H��$$  Q�����o�~P(�f�f/�vf(�f/�vf(�fn���M����Y��XD$�D$��4� �  �Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn�4�����Y��XL$�L$��   ���� t^�Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn����M����Y��XD$�D$��� tL�Q�L$<Q�t$�@H��$�   Q�����o�~P(�f�f/�vf(�f/�vf(�fn���+����L$�E���M�T$$��D$(@�D$(���T����t$,�EF�t$,�X������fW`�f(��L$�Y��L$�Y��X��L$0�Y��X��Nn ����^ȋE_^�\$�D$�d$(f�(��Y\$��$�   ��$�   ����Y��Y��Y��Y��Y��X��X��X�f��f�`��]� �U����y Vt�u�u�u�uV�q5  ��^��]� �Mj ��  ��W�WɅ�t/�D�j V�A@�@8�Ѓ��M��u�uVQ���RH�o �~H�E^� f�H��]� U���   VW��� t�u�u�u�uV��4  _��^��]� �MSj �F  ��W���u�E[_^� f�@��]� �uW��M�f�x���fE�fE�fE���tjh��x���VP�p ��WɃ4�o�~f�E�����e��e��Z  �~T �P  ��# �ȉE�
$ j���   P�� ���P�2 �M���o��M�oB�A�M�oB �A �E�oB0�@0�E�oB@�@@�E�oBP�@P�E�Oxf�@fY�@�@(�Y��@(@0���   f�fY�@0�@@�Y��@@@H���   f�fY��YHX@H�HX�E�oG`� �E�~Gpf�@�� ����uP�1h���M���o �A`�o@�Ap�o@ ���   �o@0���   �o@@���   �o@P���   �Eƀ�    �Eƀ�    �E�O4���   �E�G@���   �E�GH���   �E�GP���   �E�GX���   �Eǀ�      �Eǀ�       �Eƀ  �8 t
�E���   �< t
�E���   �M̍E�P���   P���   P�uQ�������u�o�x����E��~E�f�E��EP�! �E����E��   �oP�U��]��\W@�\_Hf.���D{�^��(��oXf.��U���D{�^��(ك8 �]�uYf/�v(��	f/�v(�f/��e�v(��	f/�v(�f/�v(��	f/�v(�f��U��e��8 ��   �< �E���   ���N �]��E����N �]�W�f/����]�v	�X��]��U�f/�v	�X��U����f/�v�\�(��\��E�f/�vY�\��\��M��J���N �]��E����N �U�W�f/�����]�v	�X��U��U�f/�v	�X��U��E�3�9��   �oE�E��E̡D���x���Q�E�f�E��@@S�@8�Ѓ���x�����uQS��`���Q���RH[_^�o �~H�E� f�H��]� ���������������U������  ��3ĉ�$�  �ES�]VW���\$(�M�|$ �D$,� t�uPQS���/  �(  �HTW�W�f(��
  ���  ;GL��  �_@f/���  �H �o��   ��$�   �~��   fք$�   u"�o��   ��$�   �~��   fք$�   �4 W���������,�f�$�  D���$�  f�$  f�$   f�$0  f�$@  f�$P  f�$`  f�$p  f�$�  f�$�  ��$  ���   �@0��$�   ��$  ( �P��$�  f֌$�  ���   ��P��$�   P�t> �T$8�\$\���o�RTS��$�   �~@��@  �D���$  fք$�  fք$�  fք$l  ��$�  Q��$x  ����$�   ��$h  �o��   ��$�   �~��   ��$�   fք$`  fք$H  fք$0  W�fD$p�D$h    f�$�   �D$d    f�$�   Ǆ$�       �$�   fn������$P  ��$8  ��$   �@�$QR��   ��$�   Q�Ѓ��o�\$(�~@�D$P�D$HfL$0���   ���\$,���@	��   ��$�   �|$P��$�   ��$   �ST�D��Y�W�Yˍ�@  Q�YӍ�$�   ���\$p�X��D$x�X���$�   �X�f�fn������$�   f֌$�   ��$P  f֌$`  ��$8  f֌$H  ��$   f֌$0  �@�$QR��   ��$�   Q�������o�~@�D$PfL$0��������|$ �\$(�D$H�G4H��   H�H  9D$T�8  �T$`�D$h�\�$�   �\�$�   �L$p�\�$�   �Y��Y��Y��X��X��c ���D$G8$�g����荄$�   �OP����\$(�D$(�$P�� ���@�$�q�|$T ��   �T$`�D$h�\�$�   �\�$�   �L$p�\�$�   �Y��Y��Y��X��X��!c ���D$G8$�����������$�L���D$8���\$ �L$ f�fY�D$0�D$H�Y�fL$0�W�W��f�C��$�  ��_^[3��G ��]� ���U���|S��V�]��{ t�u�u�u�uV�;*  ��^[��]� W�}W�fE��E�OT����  �{@ �o��   �E��~��   f�E�u�o��   �E��~��   f�EġD�Q�@�@X��3ɉE���M����  �D�Q�wT�@�@T�Ѓ����{L �u�t8�D����   �M�RT���v�KLP�K 3�9SH��3Ƀ����;��   �GT���   ��@  ���}��]����   �]���   ���   �D��{T�]��@��(  �}���p  W�}jSRQ�M�Q�OTV�u�Q�M�Q�Ћ]���,�o �{D �~X�E��C8�M��U��Y��Y��Y��X]��XM��XU�th���f(�W��e�f/�v�]��f/�v�E�f/�v(��	f/�v(�f/�v(�f��M��#f/�v(�f��M���M��U��]�MA�M;M��y����E�oE�_^� [�E�f�@��]� ����U���0VW��� t�u�u�u�uV��'  _��^��]� �Mj �J  ����u�EW�_^ �@��]� �D�j V�@@�@8�Ѓ��M��u�uVQ���RH�oE�G4�M�W�����EЃ�w&�$��<�E��E���M���]���U�G8�E��eЃ�w(�$��<�e���E���M���]���U��G<��w�$��<(��(��(��(ʋE�oE�_^� f�H��]� �/<<</<#<*<H<O<V<i<]<d<x<}<�<�<�<�<����U����   SVW���}�� t�u�u�u�uV�g&  ��_^[��]� �]W�W��{T �	  �Mj �  ( �������U�f�4�����t=�D�j V�A@�@8�Ѓ��������uSVQ���RH�o ��4����~@�E��P W��KTW�fE��M��o��   �E��~��   f�E�u�o��   �E��~��   f�E��G@3�9��  �Yx���3�9WTQD�3��E��X��D��u�@�E��@X�Ѓ�����  �E��E��E��E���I �D�V�sT�@�@T�Ћ؃��]؃�$   �n  �\ t8�D����   �M�@T���s�O\P� 3�9WX��3Ƀ����;��0  �GH�]�U��M��e��[T�Y�j �Yȍ�@  �D����   ���   �Y����   j���   �X��X�W��X��   �M��]��E�W�f�|����e�f�d�����t�����(  ���   �@��V�u��u؋�d  WRQ�M�Q�M�Q��d���Q��|���QVS�Ѓ�8���S  �}���  �E�    �E�    �9 t$�E�P�E�P�GT��0  Q�/F ���}� �  ���   ��   �D�W��WTW�f����f�L����E���,�����\����H��L���P�����P��(  ���   P�E�P�E�P���   ��P��`  ���$j jVR����L�����4��T�����\����Y�|����}��YU��Y]��G8�Y��Y��Y��XM��XU��X]��M��U��]��,  ��l�����d���f(��M�f(��e���t����U��Y��GT�Y܋��   �X�f(��Y��X��@ �Y��Y��Y��Y��\��H�\��\��Y��Y��X��H(�Y��X�W�f/���   �M��M f(�W�f(�f(��YM��Y�|����YU�f/�vf(�f/�vf(�f/�vf(؋}��G8�Y��Y��Y��E��X��E��E��X��E��E��X��E���}��D��]�E�@�sT�@X�Ћu��;��H����E��M��
�M��E��Y�4����Y�<���f(��E��YE�fыE_^[�f�@��]� �����������U��y Vt�u�u�u�uV�!  ��^]� �q4�M�b  ����u�EW�^ �@]� �D�j V�@@�@8�Ѓ��ȋ�u�uV�uV�RH��^]� �������������U����y t�u�u�u�u�   �E��]� �I4��t1�D��U��uR�@ �@X�ЋM�o ��~@��f�A��]� �EW� �@��]� ��������������U����   �y Vt�u�u�u�uV��  ��^��]� �u��SWj �W
  j�΋��L
  j�΋��A
  j�ΉE�5
  �uW��E�W��M�fE�fE�fE�fE���tjh��|���VP�[ ����E��E�����< �Fݝ|����E��E�����< �%��W�f/��|����]�v�X�f/F�U�v�X����3�3�f/ٍQrf/�G�f/�rf/�GA���m  �$�F���^  ���E��Y�W�Y��Y���|����U��E��"������|����uQW��d�����   ���  ���E��Y�S�Y��Y��\��U��E���|����B"������|����uQ������   �]����   ���E��Y�S�Y��Y��\���|����E��U���!������|����uQ��4����S�]��tc���E��Y�S�Y��Y��\��\��E���|����U��!������|����uQ��L���S�Q���RH�o fE��~@�EfM�_[�^f�@��]� ��D�D6E�EU���   VW��� t�u�u�u�uV�;  _��^��]� �G`W�� �f.����Dz�W`�Ghf.����Dz�Wh�Mj �d  ����u�EW�_^ �@��]� �EW��G8�%`�f.��o��U��]��\Wp�\_x�U��]���D{	fW��U��G@f.����D{	fW��]��GX��R �E��GX��B �oe���`���f(��E�f(�f(��YU�jh�YE��Y��Y��\��X��^_`�^Wh�\_H�XWP�X_p�XWx�}WP�]��U��W �oM�D��E�f��~G��`���j fօp����@@V�@8�Ѓ���`�����uQV�u��V�RH_��^��]� ���������������U��E�A�E    ]���  ����������U��D�SV�u�ً@@WV�@,�ЋD����΋����   �RT�ҋD�j Ph�  �Q�ϋBl�ЋD���j h�  �Q�ϋ��   �ҋ���u
_�s^[]� �D��΋��   �@��=�� u
_�s^[]� �D��΋��   �@��=�� t�D��΋��   �@��=�� u���  P�:�������P��  �C_^[]� �����U��W�f/Ev����E�E]�����E�E]����������������U���X�D��M�SVQ�@�@�СD��M�j j�h���@Q�@�СD��M�E�    ���@�@<�ЋD��؍E�P�I�I�ыD�j j�h���A�M�Q�@�СD��M����@j�Q�M�@DQ�M�ЋD����E�P�I�I�у�����  W�}��C�;�u}�D��M�Wj Q�@�M�@P�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��MQ�M�Q�@�@�СD��M�Q�@�@�Ѓ��-  G;��$  ��$    �D��M�jWQ�@�M�@P�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M����E�    �@j Q�M�@@Q�M��Ѕ��D��@��   �u��@P�M�j Q�M�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��MQ�M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@��G�� ;��������@�M�Q�Ѓ�_�D��uV�@�@�СD��MVQ�@�@�СD��H�E�P�I�ыD��EP�I�I�у���^[��]� ���������������V���L  �����  j jjZjZ�ȉF0�ۈ  �N0j j j 轉  �F    ���F   �F    �F   �F   �F    �F    �F$   �F(   �F,    ^����VW��j j h,� �����h �O0�w0��蚇  V脋  ����_^�L  ��������U��D�SV���   �@(�Ћ]����t\W��tT�D�V�@@�@,�ЋD��������   �΋RT�ҋD�h*� Ph�� �Q�ϋBl��;�tj ����������u�3�_^[]� _��^[]� �������U��D�SV���   �@,�Ћ]����t\W��tT�D�V�@@�@,�ЋD��������   �΋RT�ҋD�h*� Ph�� �Q�ϋBl��;�tj ����������u�3�_^[]� _��^[]� �������U��D�V��W�@@V�@,�ЋD����΋����   �RT�ҋD�j PkEd�Q���� P�Bl��_^]� �D����   �@x��U��} �   V�   E�D�Q�@@�@��#�3Ƀ�;�����^]� ���������̡D�V��V�@@�@�Ѓ��u�D�V�@@�@�Ѓ��u3�^ø   ^��������̡D�V��W�@@V�@,�ЋD����΋����   �RT�ҋD�h*� Ph�� �Q�ϋBl��_^���������U���0�D�Q�@@�@,�ЋD���W���fE��E��A�M�Qh�� �MЋ��   Q�����o�~@�Ef�E���Ef����]� ����U���0�D�Q�@@�@,�ЋD���W���fE��E��A�M�Qh�� �MЋ��   Q�����o�~@�Ef�E��f��H��]� �����̡D�Q�@@�@,�ЋD����ЋA��j h=  ���   �����U��D��� �@@VWQ�@,�ЋD����E�P�I�I�ыD����A�M�Qh;  �M����   Q���ЋD����}W�I�I�ыD�WV�A�@�СD��H�E�P�I�ыD��E�P�I�I�у���_^��]� ���������������U��D��� �@@VWQ�@,�ЋD����E�P�I�I�ыD����A�M�Qh<  �M����   Q���ЋD����}W�I�I�ыD�WV�A�@�СD��H�E�P�I�ыD��E�P�I�I�у���_^��]� ��������������̡D�Q�@@�@,�ЋD����ЋA��j h>  ���   �����U��D��� �@@VWQ�@,�ЋD����E�P�I�I�ыD����A�M�Qh?  �M����   Q���ЋD����}W�I�I�ыD�WV�A�@�СD��H�E�P�I�ыD��E�P�I�I�у���_^��]� ��������������̡D�V�񋀈   �@T��j P���u  ^��U��D�VW���@@W�@,�ЋD���kMd���B�u���� Q�@p���Ѓ} tjW���  j j h,� �b ��_^]� �U��D����   �@|]��������������U��} �   SVW�   ��E��D��} Stw�@@�@��#ǃ�;�t�D�S�p@�F���P�FS�Ѓ��} t\�D��ˋ��   �@P�Ћ���tD�D����   �ˋRL�ҋD�S���   �΋@h��_^[]� �p@�F����#�P�FS�Ѓ�_^[]� �������U��D�Q�@@�@,�ЋD����ЋA���uh�� �@p��]� ��������������U����D�Q�@@�@,���E���D����E��E�E�W��E��A�M�Qh�� �ʋ@H�Ћ�]� ������������U����D�Q�@@�@,��E�D�����E�W��E��A�M�Qh�� �ʋ@H�Ћ�]� ��������U��D�V��V�@@�@,�ЋD����ȋB�uh=  �@0��jV���w  j j h,� �y` ��^]� �U��D�Q�@@�@,�ЋD����ЋA���uh;  �@8��]� ��������������U��D�W��W�@@�@,�ЋD����ȋB�uh>  �@0�Ѓ} t
j W����  j j h,� ��_ ��_]� �����������U��D�Q�@@�@,�ЋD����ЋA���uh?  �@8��]� �������������̡D�VW���@@W�@,�ЋD������΋Rj h=  ���   �ҋD��Q3Ʌ����B0Qh=  ����jW���(  j j h,� �*_ ��_^����̡D�SV�ً@@WS�@,�ЋD������ϋRj h>  ���   �ҋD����Q3Ʌ����R0Qh>  ���҅�u	VS���   j j h,� �^ ��_^[��������������U��D�Q�@@�@�ЋЃ�#U3�;U��]� �����������U��D�VW���p@W�F��EP�FW�Ѓ�_^]� ��������U��D�VW���p@W�F�ЋU��#�P�FW�Ѓ�_^]� ����U��D���4�@SV�ٍM̋@WQ�СD��\��u��j j��H�T�D�P�E�P�A�СD��M�Q�@�@�СD��M�j j�hd��@Q�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M��4�@�@<�ЋD�j�j��Q�M�QP�M�BL�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��}W�@@�@,�ЋD����ЋA��jh�  �@0�СD��ϋ��   �@��-�� �Q  ���@  ��&�7  ���7  �D��ϋ��   �@P�ЋD��Ћ��   �ʋ@X�Ћ؅��  ��    �D�j S�A@�@8�Ћȃ�3��M��E��� �P�R\��tZ�D�S�@@�@,�ЋD��������   �ˋRT�ҋD�j PV�Q�ϋBl�Ћ};�u�D���j hȴ ���   �@�ЋE��d�M�@�E��Q� |��D�W�@@�@,�ЋD��������   �ϋRT�ҋD�h*� Ph�� �Q�΋Bl��P��������؅�����_^[��]� W���   _^[��]� �������U��V�O �D����u�I@�I,�у���Vh�  �i  �Ѕ���   �D����   �ʋ��   �Ћ�����   W���$    �D��΋��   �@��=.� ug�D�V�@@�@,�ЋD������Q��j h�  ���   �ҋD��P3���?B OЋARh�  �ϋ@4�СD���j j���   �@�СD��΋��   �@(�Ћ����d���_^]� ��������������U����D�V�uV�@@�@,�ЋD�W����E���fE�A�M�Qh�� �ʋ@H�СD�V�@@�@,�ЋD������Q��j h�  �R0�ҋD�jh�  �A�΋@0�СD���j h�  �@�@4�СD���jh5  �@�@0�СD���jh6  �@�@0�СD���jh7  �@�@0�СD���j h8  �@�@0�СD���j h:  �@�@0�СD���jh9  �@�@4�СD��M�Q�@�@�СD��M�j j�h���@Q�@�СD��M����@Qh;  �΋@8�СD��M�Q�@�@�СD����΋@j h=  �@0�и   ^��]� ������U��]�go  �������U��]�p  �������U��Q�D�S�u�M��@@�@,�ЋM����j �� ���������w �D���j h8  �@���   ��[��]� �u�M��u�u�u�u�o  [��]� ��������������U����D�SVW�@@�ً}j W�@8�Ћu���E���*  t��tA���O  ���F  �D���j hȴ ���   �@��j j h,� �W ���  �M�	�E �D��M�Q�@�@�СD��M�j j�h0��@Q�@�СD��M�Q�@�@�ЋE���j Wj*�E �D��M�Q�@�@�СD��M�j j�h<��@Q�@�СD��M�Q�@�@�ЋE����'E �D��M�Q�@�@�СD��M�j j�hH��@Q�@�СD��M�Q�@�@�Ѓ��5��-�� t��u'jW��������D��ϋ��   �@T�ЋMP��Rh�u��VW�em  _^[��]� ������������U����D�S�]V���   �M���W�@�Ћ}=�� �D���   ���   �ϋ@T�Ћ��HJ ;�ug�D��M�Q�@�@�СD��M�j j�h ��@Q�@�СD��M�Q�@�@�Ћu�����j W������D���j h�� ���   �@����u��u���uWS�u�l  _^[��]� �@@W�@,�ЋD����؋��   �ϋ��   �ҋЅ�tH�D��uj ���   �ʋ �ЋD���j V�ϋ��   ���   �ҋD�Vh�  �A�ˋ@p��_^�   [��]� ���������������U��Q�D�SVW�@@�}j W�@8�Ѓ��E�3۾�� ���S�R\��tj�D�W�@@�@,�ЋD��������   �M�RT�ҋD�j PV�Q�ϋBl�Ћ���t&�D�j W�I@�I8�у��ȋ�u�uW�RD��u�}��dC��Q� }�E��v���3�_^[��]� ����U��Q�D�SVW�@@�}j W�@8�Ѓ��E�3۾�� ���S�R\��t`�D�W�@@�@,�ЋD��������   �M�RT�ҋD�j PV�Q�ϋBl�Ћ���t�D�j W�I@�I8�у��ȋW�RL�}�E���dC��Q� |�_^[��]� �����U��V�u�u���uV�{������u  �D�SWj �@@V�@8�ЋD���V�I@�I,�ыD������Q��j h�  ���   �҅��'  �D���jh�  �@�@0�СD���j h=  �@���   �ЉC�ϡD�jh�  �@���   �ЉC�ϡD�j h�  �@���   �ЉC�ϡD�jh9  �@���   �ЉC�ϡD�jh8  �@���   �ЉC�ϡD�j h:  �@���   �ЉC�ϡD�jh5  �@���   �ЉC �ϡD�jh6  �@���   �ЉC$�ϡD�jh7  �@���   �ЉC(�D����   �@T���ЉC,_3�[^]� ���������U��D�VW�}�@@j W�@8�Ѓ��ȋ�Rd��~r�D�W�@@�@,�ЋD����ϋ����   �RT�ҋD�j Ph�� �Q�΋Bl�Ћ���t.�D�j V�I@�I8�у��ȋ�u�uV�uV�RH_��^]� �EW�_^ �@]� ����U��V�u��V������D�V�@@�@,�ЋD������Q��j h�  ���   �҅�t�D���j h�  �@�@0��^]� �����U���@V�  (���M����E�fE�P�H��E���,���D��M�Q���   �@@�ЋD����Q��Ph�  �E�P���   �ЋD��u�o ���   ��~@�E��	Pf�F�у���^��]� ���̸   �����������U��D�V�uV�@�@�Ѓ}c�D�j j��I�Iuh�V�у���^]� hL�V�у���^]� ̸   � ��������U��MW��E�A��c��   ��Xf�$�Df(��������f�I]� (��������f�I]� (��������f�I]� (���X��f�I��]� ��e�ef%f=f ����3���������������U����   SVW�}���u�B ���^�]����  �N0����  �D�Q�@�@�Ѓ�����  ���k������q  �D�S�@@�@,�ЋD����؋Q��j h�  ���   �҅��<  �D���j h�  �@�@0�ЋN0��l  �N0j jjZjZ�m  �N0j j j �bn  W������WfE��E��  ������jQ�u���PD����  ������  �x�W��E�3��E�    f�E�fE��E�   ��x�������]�f�E��fn�3�����^��M����$    �d$ fnÍ�`�������jQ�M��u�^�Q��f���`���W�fօp����PH���W��of/�f]��~Pv�M��f/�v�E���]��]�f/�v�M��f/�v�E���]�f/�v(��	f/�v(��oE�D��M�f�U��E�j�@Q�M�Q���  ������ofM��~@�D��E��YH�,�(�f�P�Y��Y��,�P�,�P��  WS�v0���M�C�x���$��Z�����G��Z���������u�PL��$����4  _^[��]� ���������U��D�j �u�@@�@8�Ѓ�]�������U��E���   ����V��i�|  ���l�$�|l�E^�    �@   ��]ËE^�    �@   ��]ËE^�    �@   ��]ËE^�    �@�   ��]ËE^�    �@    ��]ËE^�    �@x   ��]ËE^�    �@   ��]ËE^�    �@
   ��]ËE^�    �@    ��]�(���EЋMfE�P����E��&���E^��]�(p���p����Mf�p���P����E��&���E^��]�( ��E��MfE�PW��E��Z&���E^��]�(����@����Mf�@���P�����P����$&���E^��]�(���E�MfE�P����E���%���E^��]�(��E��MfE�P�P��E���%���E^��]�(@��E��MfE�P����E��%���E^��]�(����X����Mf�X���P�H���h����g%���E^��]�(����(����Mf�(���P�p���8����1%���E^��]ËE^�     �@    ��]��ij#j8jMjbjwj�j�jk�j�j>ktk�k�k�k1lgl  	
��������������U���\V��I �D���h&� �A�ʋ@T�Ћ�����  �M���T  ���I �D���Vh&� �A�ʋ@D�ЍM��U  �oI �D���h&� �A�ʋ@T�Ћ���u^��]áD��M��E�   �E�   Q���   �@8�ЋD����Q��PhM  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��PhR  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��RhN  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����QP�B4��hO  �СD��M�Q���   � �СD��M��E�   �E��   Q���   �@8�ЋD����Q��PhP  �B4�СD��M�Q���   � �СD��M��E�   �E�    Q���   �@8�ЋD����Q��PhQ  �B4�СD��M�Q���   � �СD��M��E�   �E�x   Q���   �@8�ЋD����Q��PhS  �B4�СD��M�Q���   � �СD��M��E�   �E�   ���   �@8Q�ЋD�����ҋA��Rh]  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��PhT  �B4�СD��M�Q���   � �СD��M��E�   �E�
   Q���   �@8�ЋD����Q��PhU  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��Rh\  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��Ph_  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��RhZ  �΋@0�СD��M�Q���   � �СD��M��E�   �E�    Q���   �@8�ЋD�����ҋA��Rh[  �΋@0�СD��M�Q���   � �Ѓ�(���E�fE��M����P�E��C���D��M�Q���   �@@�ЋD����Q��Ph^  �BH�СD��M�Q���   � ��(p��E����M�fE����P�E������D��M�Q���   �@@�ЋD����Q��PhW  �BH�СD��M�Q���   � ��( ��E����M�fE�W�P�E��x���D��M�Q���   �@@�ЋD����Q��PhX  �BH�СD����   �M�Q� �СD��M��E�   �E�   Q���   �@8�Ѓ��M�fn��D����QhY  ��f�E��E��@�@H�СD��M�Q���   � ��(���E����M�fE����P�E�����D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE����P�E��C���D��M�Q���   �@@�ЋD����QP�BH��h�  �СD��M�Q���   � ��(��E����M�fE��P�P�E������D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(@��E����M�fE����P�E��s���D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE��H�P�E�����D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE��p�P�E�����D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � �Ѓ���^��]����������U��D��MQ�@�@�Ѓ�]��������U��V��W��F�N����F��&  �u���c�  ��^]� ������������U��VW��j j h,� �����> �O0�w0���]  V�qa  �����"  �Et	W�[$  ����_^]� U����Af.���E����Dz���]���u���]���̡D����   �@(��D����   �@,��D����   �@x��D�Q�@@�@�����������������U���0�D�Q�@@�@,�ЋD���W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�Ef�E���Ef����]� ����U���0�D�Q�@@�@,�ЋD���W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�Ef�E��f��H��]� �����̡D�Q�@@�@,�ЋD������Q�$�A��h�  ���   ������������U���0�D�Q�@@�@,�ЋD���W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�E�,�fɉ�E�,�f�E����]� U���0�D�Q�@@�@,�ЋD���W���fE��E��A�M�Qh�  �MЋ��   Q�����o�~@�Ef�E��f��H��]� ������U��D�Q�@@�@,�ЋD��Ѓ��A�Mj ���   �����  ��Q����]� �U��D����   �@|]��������������U��D�VW���p@W�F�Ѓ} t������P�FW�Ѓ�j j h�� �u; ��_^]� ������������U����D�Q�@@�@,��fnE���D�������E�fnE����E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ����U����D�Q�@@�@,��E�D�����E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ��������U��D�Q�@@�@,�ЋD����EQ�$�A��h�  �@,��]� ���������U����D�Q�@@�@,��fnE���D�������E�fnE����E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ����U����D�Q�@@�@,��E�D�����E�W��E��A�M�Qh�  �ʋ@H�Ћ�]� ��������U����D�VWQ�@@�@,�ЋD����u���A�Nd�����@0j Q���СD��4�W���fE��E��P�E�P���  P�BH�СD�������ϋP���  �$P�B,��_^��]� ������������U��D���P�@@VWQ�@,�ЋD����u���A�Nd�������   j Q���Ѕ���   �D��4�W���fE��E��P�E�P���  P�E�P���   �Ѓ����o �E��~@�D�f�E�����$�P���  P���   �СD����]��E��ϋ@�$h�  �@,�СD��M�Qh�  �ϋ@�@H��_^��]� ��������U���P�D�VWQ�@@�@,�ЋD���W���fE��E��A�M�Qh�  �M����   Q���Ѓ����o �E��~@�D�f�E�����$�@h�  ���   �СD��ϋuj�]��P�Fd����P�B0�СD��4��ϋP�E�P���  P�BH�СD����E��ϋP���  �$P�B,��_^��]� ��̸   � ��������� �������������U��E���   ����V��i�|  ��h��$���E^�    �@   ��]ËE^�    �@   ��]ËE^�    �@   ��]ËE^�    �@�   ��]ËE^�    �@    ��]ËE^�    �@x   ��]ËE^�    �@   ��]ËE^�    �@
   ��]ËE^�    �@    ��]�(���EЋMfE�P����E�����E^��]�(p���p����Mf�p���P����E������E^��]�( ��E��MfE�PW��E�����E^��]�(����@����Mf�@���P�����P�������E^��]�(���E�MfE�P����E��W���E^��]�(��E��MfE�P�P��E��*���E^��]�(@��E��MfE�P����E������E^��]�(����X����Mf�X���P�H���h��������E^��]�(����(����Mf�(���P�p���8�������E^��]ËE^�     �@    ��]Ù~�~�~�~�~,��AV��A�n���р�  	
��������������U���\V�$5 �D���h&� �A�ʋ@T�Ћ�����  �M��+@  ����4 �D���Vh&� �A�ʋ@D�ЍM��d@  ��4 �D���h&� �A�ʋ@T�Ћ���u^��]áD��M��E�   �E�   Q���   �@8�ЋD����Q��PhM  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��PhR  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��RhN  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����QP�B4��hO  �СD��M�Q���   � �СD��M��E�   �E��   Q���   �@8�ЋD����Q��PhP  �B4�СD��M�Q���   � �СD��M��E�   �E�    Q���   �@8�ЋD����Q��PhQ  �B4�СD��M�Q���   � �СD��M��E�   �E�x   Q���   �@8�ЋD����Q��PhS  �B4�СD��M�Q���   � �СD��M��E�   �E�   ���   �@8Q�ЋD�����ҋA��Rh]  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��PhT  �B4�СD��M�Q���   � �СD��M��E�   �E�
   Q���   �@8�ЋD����Q��PhU  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��Rh\  �΋@0�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD����Q��Ph_  �B4�СD��M�Q���   � �СD��M��E�   �E�   Q���   �@8�ЋD�����ҋA��RhZ  �΋@0�СD��M�Q���   � �СD��M��E�   �E�    Q���   �@8�ЋD�����ҋA��Rh[  �΋@0�СD��M�Q���   � �Ѓ�(���E�fE��M����P�E��
���D��M�Q���   �@@�ЋD����Q��Ph^  �BH�СD��M�Q���   � ��(p��E����M�fE����P�E��;
���D��M�Q���   �@@�ЋD����Q��PhW  �BH�СD��M�Q���   � ��( ��E����M�fE�W�P�E���	���D��M�Q���   �@@�ЋD����Q��PhX  �BH�СD����   �M�Q� �СD��M��E�   �E�   Q���   �@8�Ѓ��M�fn��D����QhY  ��f�E��E��@�@H�СD��M�Q���   � ��(���E����M�fE����P�E��	���D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE����P�E�����D��M�Q���   �@@�ЋD����QP�BH��h�  �СD��M�Q���   � ��(��E����M�fE��P�P�E��;���D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(@��E����M�fE����P�E������D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE��H�P�E��k���D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � ��(���E����M�fE��p�P�E�����D��M�Q���   �@@�ЋD����Q��Ph�  �BH�СD��M�Q���   � �Ѓ���^��]����������U����M�������E���u��]� SV�u��Wj 薓 j �΋�苓 �u��؍E�V�u�7P�G����M���P�3�� �D��M�Q���   � �Ѓ��   _^[��]� �����U���V��M�hM  �:� ��M�j Q���PD�M��5� hR  �M��� ��M�j Q���PD�M��� hN  �M���� ��M�j Q���PD�M��� hO  �M��ԏ ��M�j Q���PD�M��ϑ hP  �M�貏 ��M�j Q���PD�M�譑 hQ  �M�萏 ��M�j Q���PD�M�苑 hS  �M��n� ��M�j Q���PD�M��i� h]  �M��L� ��M�j Q���PD�M��G� hT  �M��*� ��M�j Q���PD�M��%� hU  �M��� ��M�j Q���PD�M��� h\  �M��� ��M�j Q���PD�M��� h_  �M��Ď ��M�j Q���PD�M�运 hZ  �M�袎 ��M�j Q���PD�M�蝐 h[  �M�耎 ��M�j Q���PD�M��{� h^  �M��^� �j �M�Q���PD�M��Y� hW  �M��<� ��M�j Q���PD�M��7� hX  �M��� ��M�j Q���PD�M��� hY  �M���� ��M�j Q���PD�M��� h�  �M��֍ ��M�j Q���PD�M��я h�  �M�贍 ��M�j Q���PD�M�诏 h�  �M�蒍 ��M�j Q���PD�M�荏 h�  �M��p� ��M�j Q���PD�M��k� h�  �M��N� ��M�j Q���PD�M��I� h�  �M��,� ��M�j Q���PD�M��'� �   ^��]� �����������U����D�S�M��M�W�@Q�@�СD��M�j j�hX��@Q�@�Ћ}�E����P蹕 ���M�D�Q�Ë@�@�Ѓ���t
_3�[��]� V�u� �  hM  �M��x� �]��M�WQ�ˋ�PD�M��q� hR  �M��T� ��M�WQ���PD�M��P� hN  �M��3� ��M�WQ���PD�M��/� hO  �M��� ��M�WQ���PD�M��� hP  �M��� ��M�WQ���PD�M��� hQ  �M��Ћ ��M�WQ���PD�M��̍ hS  �M�诋 ��M�WQ���PD�M�諍 h]  �M�莋 ��M�WQ���PD�M�芍 hT  �M��m� ��M�WQ���PD�M��i� hU  �M��L� ��M�WQ���PD�M��H� h\  �M��+� ��M�WQ���PD�M��'� h_  �M��
� ��M�WQ���PD�M��� hZ  �M��� ��M�WQ���PD�M��� h[  �M��Ȋ ��M�WQ���PD�M��Č h^  �M�觊 ��M�WQ���PD�M�裌 hW  �M�膊 ��M�WQ���PD�M�肌 hX  �M��e� ��M�WQ���PD�M��a� hY  �M��D� ��M�WQ���PD�M��@� h�  �M��#� ��M�WQ���PD�M��� h�  �M��� ��M�WQ���PD�M���� h�  �M��� ��M�WQ���PD�M��݋ h�  �M���� ��M�WQ���PD�M�輋 h�  �M�蟉 ��M�WQ���PD�M�蛋 h�  �M��~� ��M�WQ���PD�M��z� ��]����VW�u�f:  ^_[��]� �������������U���   SVW���]����}�؅��/  j ���� ���������i�  ����$�ܔj ���ߋ �0�E�P�����D�P���   �@8�Ѓ��ϋ�j 贋 �D�V�0�Q�ˋ��   �ЉE�M�D��E�   j Q���   �u�@�СD��M�Q���   � �ЍM��D�Q���   � �ЋE����   _^[��]� j ���5� �0�E�P����������p���j �ϋ��� �D�V�0�Q�ˋ��   �ЉE؍MСD��E�   j Q���   �u�@�СD��M�Q���   � �ЍM��\���j ��踊 �0�E�P�}����D�P���   �@@�Ѓ��ϋ�j 荊 �D�V�0�Q��p���P�ˋ��   �ЍM�Q�M��o Q�E��~@�D�f�E��E�    �E�    ���   �@�СD��M�j Q�u���   �@�СD��M�Q���   � �СD��M�Q���   � �ЋE����   _^[��]� �u���uW�u� 8  _^[��]� �I ��b�ߓ��          ����������U��SVW���s����}�؅���  j ���� ���������i�~  ��H��$�,��D��u���   �@8�Ѓ��ϋ�j �݈ �D�V�0�Q�ˋB4�ЋE_^[��   ]� �D��u���   �@8�Ѓ��ϋ�j 藈 �D�V�0�Q�ˋB0�ЋE_^[��   ]� �M�����j �ϋ��_� �D�V�0�Q�B0����j j h,� �E�� ���   _^[]� �D��u���   �@8�Ѓ��ϋ�j �� �D�V�0�Q�B4맡D��u���   �@@�Ѓ��ϋ�j �և �D�V�0�Q�BH�r����M����j �ϋ�诇 �D�V�0�Q�ˋBH��j j h˴ �K����u���uW�u��5  _^[]� �����w���.�ޖ�  ��������������U��D�Q���   �@X�Ћȃ���u]� �D��u�u�@|Q�@�Ѓ�]� ����U��D�Q���   �@X�Ћȃ���u]� �D��u�u�@|Q�@8�Ѓ�]� ����U��UV��j j j ��D�R�@�@�Ѓ��F��^]� ���̡D�Vj ��@j j �6�@�Ѓ��F^�U��V��N��u3�^]� �D�Q�u�@�u�6�@�Ѓ��F�   ^]� �����������������������������̅�t�j������̡D��@��  ��D��@��(  ��U��D��U���@R��   �ЋMP�  �M���  �E��]� �����������̡D��@��$  ��U��D��@��  ]��������������U��D��@���  ]�������������̡D��@��  ��U��D��@���  ]��������������U��D��@��x  ]��������������U��D��@��|  ]�������������̡D��@��d  ��U��D��@��p  ]��������������U��D��@��t  ]��������������U���EV����t	V�   ����^]� ��������������U��D��E��t;�} �   �u�I�ut;�B�P���   �Ѓ�]Ã�B�P���  �Ѓ�]ù   ;�VB�W�xW� ������u_^]À} tWj V�D
 ��������F_���   ^]�����������U��M��t+�=�� t�y���A�u	�E]�� �D��@�M� ]��]����������U��M��t�D��@�M��@  ]��]áD�hﾭދ@��@  ��Y����������U��V�u���t�D�Q�@� �Ѓ��    ^]�����������U��D��@���  ]��������������U��E��t�x��u�   ]�3�]������U��D��@��  ]�������������̡D��@��   ��U��E�   ;�VB�W�xW� ������u_^]Ã} tWj V�� ��������F_���   ^]���������������������������������������������������������������̡D��@$�@X�����U��D��@$�@\]�����������������U��D��u�u�@$�uQ�@`�Ѓ�]� ��������������̡D�V��V�@�@�СD�V�@$�@D�Ѓ���^�����������U��D�V��V�@�@�СD�V�@$�@D�СD��uV�@$�@d�Ѓ���^]� ���U��D�V��V�@�@�СD�V�@$�@D�СD��uV�@$�@�Ѓ���^]� ���U��D�V��V�@�@�СD�V�@$�@D�СD�V�u�@$�@L�Ѓ���^]� ��̡D�V��V�@$�@H�СD�V�@�@�Ѓ�^�������������U��D��uQ�@$�@L�Ѓ�]� �����U��D��@$�@]����������������̡D�Q�@$�@�Ѓ����������������U��D����@$VWQ�@�M�Q�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]� ���U��D��uQ�@$�@�Ѓ�]� �����U��D����@$VWQ�@ �M�Q�ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у� ��_^��]� ����U��D����@$VWQ�@$�M�Q�ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у� ��_^��]� ����U���,�E�VWP�o����D�P�E�P�I$�A�ЋD����}W�I�I�ыD�WV�A�@�СD��M�Q�@�@�СD��H$�E�P�IH�ыD��E�P�I�I�у� ��_^��]� ������̡D�Q�@$�@(��YáD�Q�@$�@h��Y�U��D��uQ�@$�@,�Ѓ�]� �����U��D��uQ�@$�@0�Ѓ�]� �����U��D��uQ�@$�@4�Ѓ�]� �����U��D��uQ�@$�@8�Ѓ�]� �����U��D��u�u�@$Q�@P�Ѓ�]� ��U��D��uQ�@$�@T�Ѓ�]� �����U��D��@$�@l]����������������̡D��@$�@p�����U��D�V��V�@$�u�@L�Ѓ���^]� ���������������U��D�V�uV�@�@�СD�V�@$�@D�СD�V�u�@$�@L�ЋD��uV�I$�I@�у���^]���U��D�V�u��@$V�@@�Ѓ���^]� ���������������U��D��uQ�@$�@<�Ѓ�]� �����U��D��uQ�@$�@<�Ѓ����@]� U��D����@$VWQ�@t�M�Q�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]� ���U��D��@(�@]����������������̡D��@(�@�����U��D��@(�@]�����������������U��D��@(�@]�����������������U��D��@(�@ ]�����������������U��D�j�u�@(�u�@��]� ����U��D��u�u�@(�u�@$��]� ��̡D��@(�@(����̡D��@(�@,����̡D��@(�@0�����U��D��@(�@4]�����������������U��D��@(�@X]�����������������U��D��@(�@\]�����������������U��D��@(�@`]�����������������U��D��@(�@d]�����������������U��D��@(�@h]�����������������U��D��@(�@l]�����������������U��D��@(�@p]�����������������U��D��@(�@t]�����������������U��D��@(�@x]�����������������U��D��@(���   ]��������������U��D����@V��M�Q�@�Ѓ��E���P�   ��u3���D��M�Q�u�@$�@�Ѓ��   �D��E�P�I�I�у���^��]� ������U��Q�D��U�R�@(�@X�Ѕ�u��]� �E3�8M�����   ��]� ���������U����D��E�    �E�    V�@(��M�Q�΋@h�Ѕ�t�M��D���u@�@�M�Q�@�СD��M��uQ�@�@�СD��M�Q�@�@�Ѓ��   ^��]� �@h@�hj  Q���   �Ћȃ��D��M��@(��u�@4��j���3�^��]� �@j �u�Q���Ѕ�u�E�P������3�^��]� �D�j �H�E�HP�u��A�u�ЍE�P�q������   ^��]� ��U��D�VW�}��@(W�@p�Ѕ�t9�D��΋P(�GP�Bp�Ѕ�t"�D��΋P(�GP�Bp�Ѕ�t_�   ^]� _3�^]� ���U��D�VW�}��@(W�@t�Ѕ�t9�D��΋P(�GP�Bt�Ѕ�t"�D��΋P(�GP�Bt�Ѕ�t_�   ^]� _3�^]� ���U��D�SVW�@(��}W�@p�Ѕ���   �D��΋P(�GP�Bp�Ѕ���   �D��΋P(�GP�Bp�Ѕ�to�D��_S�΋@(�@p�Ѕ�tX�D��΋P(�CP�Bp�Ѕ�tA�D��΋P(�CP�Bp�Ѕ�t*�G��P������t�G$��P������t_^�   []� _^3�[]� �����U��D�SVW�@(��}W�@t�Ѕ���   �D��΋P(�GP�Bt�Ѕ���   �D��΋P(�GP�Bt�Ѕ�to�D��_S�΋@(�@t�Ѕ�tX�D��΋P(�CP�Bt�Ѕ�tA�D��΋P(�CP�Bt�Ѕ�t*�G0��P�-�����t�GH��P������t_^�   []� _^3�[]� �����U��D��@(�@8]�����������������U��D��@(�@<]�����������������U��D��@(�@@]�����������������U��D��@(�@D]�����������������U��D��@(�@H]�����������������U��D��@(�@L]�����������������U��D��EQ�$�@(�@P��]� �U��D����E�@(�$�@T��]� ���������������U��D��u�u�@(�@|��]� ������U��D��u�u�@(���   ��]� ���U��D��� �@$VW�u�@���M�Q�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�Ѓ��E���P�L   �D����E�P�I�I�у���_^��]� �����������U��D��} �P(�����E�B8]����U��Q�D�VW���M�@j �@d�ЋD�h@�h�  �p�IV���   �ыȃ��D��M���u�@(��j��@4��_3�^��]� �@j VQ�M�@h�СD���V�@(�@H�Ѕ�t�D���V�u��@(�@ �Ѕ�t�   �3��E�P�T�������_^��]� �������U��D�VW�}��@(Q��@P�$�Ѕ�tG�D��GQ���$�@(�@P�Ѕ�t)�D��GQ���$�@(�@P�Ѕ�t_�   ^]� _3�^]� ������������U��D�VW�}���@(����@T�$�Ѕ�tK�D����G�΋@(�$�@T�Ѕ�t+�D����G�΋@(�$�@T�Ѕ�t_�   ^]� _3�^]� ������U��D�VW�}��@(Q��@P�$�Ѕ���   �D��GQ���$�@(�@P�Ѕ���   �D��GQ���$�@(�@P�Ѕ���   �D��GQ���$�@(�@P�Ѕ�te�D��GQ���$�@(�@P�Ѕ�tG�D��GQ���$�@(�@P�Ѕ�t)�G��P�.�����t�G$��P������t_�   ^]� _3�^]� ��������U��D�VW�}���@(����@T�$�Ѕ���   �D����G�΋@(�$�@T�Ѕ���   �D����G�΋@(�$�@T�Ѕ���   �D����G�΋@(�$�@T�Ѕ�ti�D����G �΋@(�$�@T�Ѕ�tI�D����G(�΋@(�$�@T�Ѕ�t)�G0��P������t�GH��P������t_�   ^]� _3�^]� �����������̡D��@(� ������U��D�V�u�@(�6�@�Ѓ��    ^]���������������U��D��@(���   ]��������������U��D��@(�@]����������������̡D��@(�@�����U��D�V�u�@(�6�@�Ѓ��    ^]���������������U��D��u�u�@,Q�@�Ѓ�]� �̡D��@,�@����̡D��@,�@����̡D��@,�@����̡D��@,�@ ����̡D��@,�@(����̡D��@,�@$�����U��D��@,�@]�����������������U��D��U���@,VWR�@�ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у���_^��]� ����̡D�j j �@,� �Ѓ��������������U��D�V�u�@,�6�@�Ѓ��    ^]��������������̡D��@,�@4����̡D��@,�@8�����U��D��U���@,VWR�@<�ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у���_^��]� �����U��D��U����@,VW�u�@@R�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]� ̡D��@,�@,�����U��D�V�u�@,�6�@0�Ѓ��    ^]���������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��u�u�@�@\��]� ������U��D��u�u�@��  ��]� ���U��D����E�@�$�@ ��]� ���������������U��D��EQ�$�@�@$��]� �U��D����E�@�$�@(��]� ���������������U��D��@�@,]�����������������U��D��@�@0]�����������������U��D��@�@4]�����������������U��D��@�@8]�����������������U��D��@�@<]�����������������U��D��@�@@]�����������������U��D��@�@D]�����������������U��D��@�@H]�����������������U��D��@�@L]�����������������U��D��@�@P]�����������������U��D��@���   ]��������������U��D��uQ�@��  �Ѓ�]� ��U��D��@�@T]�����������������U��D��@�@X]�����������������U��U��u3�]� �D�RQ�@ �@(�Ѓ��   ]� �����U��D��@���   ]��������������U��D��@�@`]�����������������U��D��@�@d]�����������������U��D��@�@h]�����������������U��D��@�@l]�����������������U��D��@�@p]�����������������U��D��@�@t]�����������������U��D��@���   ]��������������U��D��@��  ]��������������U��D��@�@x]�����������������U��D��@�@|]�����������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��uQ�@��  �Ѓ�]� ��U��D��@���   ]��������������U��D��@���   ]��������������U��U��t�D�RQ�@ �@$�Ѓ���t	�   ]� 3�]� �U��D�Q�u�@ �u�@L�Ѓ�]� ��U��D��@���   ]�������������̡D��@���   ��U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]�������������̡D��@���   ��U��D��@���   ]�������������̡D��@���   ��D��@���   ��D��@���   ��D��@���   ��D��@���   ��U��D�V�uV�@���   �Ѓ��    ^]�������������U��D��@� ]��D��@�@�����U��D��@���   ]��������������U��D��@��   ]��������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@�@]�����������������U��D��@���  ]��������������U��D��@�@]�����������������U����E�V�u��P�����D��M�Q�@$�@�Ѓ���t]�D��M�jQ�@�@�Ѓ���u�E�P��������t3�D�jV�@�@�Ѓ���u�D�V�@�@�Ѓ���t�   �3��D��H$�E�P�IH�ыD��E�P�I�I�у���^��]��������U��D��@�@ ]�����������������U��D��@�@(]�����������������U��D��@��  ]��������������U��D��@��   ]��������������U��D��@��  ]��������������U��D��@��  ]��������������U��D��M���@VWQ�@$�ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у���_^��]��������U��D��M���@VWQ���  �ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у���_^��]�����U��j�u�  �E��]������������U���<�P��E�    SVW��t�EĻ   P�h������-�D��M�Q�   �@�@�СD��M�Q�@$�@D�Ѓ��}�D��uV�@�@�СD�V�@$�@D�СD�VW�@$�@L�Ѓ���t(�D��M�Q����@$�@H�СD��M�Q�@�@�Ѓ���t&�D��H$�E�P�IH�ыD��E�P�I�I�у�_��^[��]������U��D��M���@VW�u���  Q�ЋD����}W�I�I�ыD�W�A$�@D�СD�WV�@$�@L�СD��H$�E�P�IH�ыD��E�P�I�I�у� ��_^��]��U��D��@��D  ]��������������U��D��@��H  ]��������������U��D��@��L  ]��������������U��D��M����@VW�u���  �uQ�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]��������������U��D��@���  ]��������������U��D��@���  ]�������������̡D�Vj j��@��@�Ћ�^���������U��D�Vj �u�@��@�Ћ�^]� �U��D�V�u��@j��@�Ћ�^]� ̡D��@�@�����U��D�Vj ��M�@j V���   �Ћ�^]� �����������U��D��uQ�@�@�Ѓ�]� �����U��D��uQ�@�@�Ѓ����@]� U��D�h#  �u�@�u�@l��]� �U��D�hF  �u�@�u�@l��]� �U��D��u�@�@t�ЋD�P���   �@X�Ѓ�]� ����U��D��u�@�@t�ЋD����uR���   �@`�Ѓ�]� ���������������U��D��u�@���   �Ћȅ�u]� �D�Q���   �@�Ѓ�]� ��������U��D��@���   ]���������������A    ���    �A    �A   ���U��D��u�u�@@�uQ�@�Ѓ�]� ���������������U��D��uQ�@@�@�Ѓ�]� �����U��D��u�u�@@Q�@�Ѓ�]� ��U��D��uQ�@@�@ �Ѓ�]� �����U��D����   �@]��������������U��D����   �@]��������������U��D����   �@ ]�������������̡D����   �@$��U��D����   ���   ]�����������U��D����   ��D  ]�����������U��D��uQ�@@�@L�Ѓ�]� ����̡D�Q�@@�@H�Ѓ����������������U��D����   ���   ]�����������U��D����   ���   ]����������̡D�Q�@H���   �Ѓ�������������U��V��M��t2�D��U���   ��t�@@R��^]� �U�@D��tR��^]� V��^]� �����������̡D��@@�@0�����U��V�u���t�D�Q�@@�@�Ѓ��    ^]����������U��D�V��V�@@�@�ЋЃ��E��t��#��СD�RV�@@�@�Ѓ�^]� �U���u �E�D������   �$�u�u���   �u�u��]� ����������U��D����   ���   ]����������̡D�Q�@H���   �Ѓ�������������U��D��uQ�@H��d  �Ѓ�]� �̡D��@@�@T�����U��D��@@�@X]�����������������U��D��@@�@\]����������������̡D��@@�@`�����U��D��@@�@d]�����������������U��D��@@�@h]�����������������U��D��@@�@l]�����������������U��D��@@���   ]�������������̡D��@@�@t����̡D��@@�@x�����U��D��@@�@|]����������������̡D��@@���   ��U��D��@@���   ]�������������̡D��@@���   ��D����   �@t��U��D��@@���   ]��������������U��D��@@���   ]��������������U��D��@@���   ]��������������U��D��@@���   ]��������������U��D��@@���   ]��������������U��D��@@���   ]��������������U��D��@@���   ]��������������U��V�u���t�D�Q�@@�@�Ѓ��    ^]���������̡D��@@�@0�����U��D��MjQj �@@�@4�Ѓ�]����U��D��MjQh   @�@@�@4�Ѓ�]�U��D��u�u�@@j �@4�Ѓ�]���̡D��@|� ������U��V�u���t�D�Q�@|�@�Ѓ��    ^]���������̡D��@|�@ �����U��V�u���t�D�Q�@|�@(�Ѓ��    ^]����������U��D��@ �@H]�����������������U��}qF uGW�}��t>�D����u���   �@D�СD��u�@@�@,�ЋD����ЋA��W�u�@p��_]������������U��D��@��T  ]��������������U��D�SVW�@@�u�@,�ЋD����u�I@�I,�ыD������y��h��hE  ����Ph��hE  ������P��T  �Ѓ�_^[]�����̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������3�� �����������3�� �����������U��M�E�A4�E�A �E��E�A0�E�A��A8#��A<(��A@7��AD-��AHs��ALn��AP2��Al]��AX_�A\b��A`l��Adg��ATX��AhZ�Apd�Atq��A(�A,    ]��������������U���   h�   ��`���j P�t� j �u��`����u�u�uP�����E h�   �E���`���P�u�uj��  ��8��]�����U���   V����	  �����   S�u�M��i����D��M�Q�@�@�СD��M�j j�h���@Q�@�Ѓ��E��M�P�/���j j��E�P�E�P��d���P������P�E�P�j�����P�E�P�]������P�  ���M����d����M��\�����d����Q����M��I����D��M�Q�@�@�Ѓ��M��-�����[t	V�"	  ����^��]� ������U��V�u���  �����^]� ������Q��  YË�`��`$��`0��`4��`8��`@����������3���������������U��E�     3�]� �������������̋�PP�   ����U����   V�u��u3�^��]�h�   ��@���j P�u� �E����@����΍�@�����`���ǅD����h�   P��u�E�(��E�7��E�-��E�n��E�s��PPj��  ��^��]�U��j�u��������u]Ë�]������`��`�������̡D��@��   ��U��D�V�u�@�6��$  �Ѓ��    ^]������������U��D�V��V�@�u��(  �Ѓ���^]� ������������U��D�Q�u�@��,  �Ѓ�]� ��U��D�Q�u�@��,  �Ѓ����@]� �������������U��E��t�P�3ҡD�RQ�@��8  �Ѓ�]� ������U��D��uQ�@��<  �Ѓ�]� ��U��D��u�u�@�uQ��@  �Ѓ�]� ������������U��D��u�u�@Q��D  �Ѓ�]� ���������������U��D��uQ�@��H  �Ѓ�]� ��U��D����@VW�u��L  Q�M�Q�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]� ������������̡D�Q�@��T  �Ѓ������������̡D�Q�@��P  �Ѓ�������������U��D��uQ�@��X  �Ѓ�]� ��U��D��uQ�@��l  �Ѓ�]� �̡D��@��0  ��D��@��4  ��D��@��p  ��D��@��t  ��D��@��\  ��U��D�V�u�@�6��`  �Ѓ��    ^]������������U���u�D��u�u�@�u�u��d  Q�Ѓ�]� ������U���u�D��u�u�@�u�u��h  Q�Ѓ�]� �����̡D�Q�@�@�Ѓ����������������U���u�D��u�u�@�uQ�@X�Ѓ�]� ������������U��D��uQ�@�@\�Ѓ�]� ����̡D�Q�@�@ ��Y�U��D����@Vh�  Q���   �M�Q�ЋD�P���   �@8�ЋD����E�P���   �	�у���^��]��������������U��D��@��   ]��������������U��D��u�u�@�uQ�@�Ѓ�]� ���������������U���u�D��u�u�@�uQ���   �Ѓ�]� ���������U��D��@�@$]�����������������U���u�D��u�u�@�uQ�@(�Ѓ�]� ������������U���u�D��u�u�@�uQ�@,�Ѓ�]� ������������U���u(�D��u$�u �@�u�u�@`�u�u�u�uQ�Ѓ�(]�$ �������������U��D�VW���@W�@�ЋD���W�J�I���u�D�H�u�u�Q�N�QPj �B4j W�Ѓ�(_^]� ���������������U���u �D��u�u�@�u�u�@4�u�uQ�Ѓ� ]� ���U��D��u�u�@Q�@@�Ѓ�]� ��U��D��uQ�@�@D�Ѓ�]� ����̡D�Q�@�@L�Ѓ���������������̡D�Q�@�@L�Ѓ���������������̡D�Q�@�@P�Ѓ����������������U��D��uQ�@�@T�Ѓ�]� �����U��D��uQ�@�@T�Ѓ�]� ����̡D�Q�@�@h�Ѓ����������������U��D��u�u�@Q���   �Ѓ�]� ���������������U��D����@V�u�u���   Q�M�Q�Ћuj PV�    �F    �D����   �I�ыD��E�P���   �	�у� ��^��]� ��������̡D��@� ������U��D�V�u�@�6�@�Ѓ��    ^]���������������U���u�D��u�u�@�u�u���   Q�Ѓ�]� ������U��D�V�u�@�6�@�Ѓ��    ^]���������������U��QS�]V��V�C    �D��@�@h�Ѓ����D�u"�@h��h�  ��0  �Ѓ�^3�[��]� �M��E    �@Q�MQ�u���   V�Ѓ���t�3�9u�~*W��I �E�<� �<�tj����
  ��t��F;u�|�_�EP�C������   ^[��]� ���U��QS�]V��V�C    �D��@�@h�Ѓ����D�u"�@h��h�  ��0  �Ѓ�^3�[��]� �M��E    �@Q�MQ�u���   V�Ѓ���tу} t�3�9u�~<W�E����t*�D�Q�@�@h�Ѓ���t�E��j�<��
  ��t�8F;u�|�_�EP�k������   ^[��]� �����������U��D��@��x  ]�������������̡D��@��|  ��D�Q�@���   �Ѓ�������������U��D��uQ�@���   �Ѓ�]� �̡D��@���   ��U��D�V�u�@�6���   �Ѓ��    ^]������������VW���O�$���W����G �G0�G@�GP�    �G`    �Gd    �Gh    �Gp�Gx�����G|   _^�����������V���X   �N^�������������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7�������xP t$V������j j j�pP�ˍGP�����H ���^�    �` t�D��w`�@�@�Ѓ��G`    _[�������������jh��h�   h�   �:�������t������3�����������U��V�uW�>��t���K����O����W蝾����_�    ^]�U��D�SVW�@��W��   �_dS�wx�w`�uV�Ѓ��G|����   �? ��   �; ��   �wpV�_hS�u���  ����u&�W���D�h��h  �@��0  �Ѓ��u�O�������跻���xP u����"��襻��j j j�pP�ˍGP葻���H ��ЉG|��t���[����G|_^[]� �G|�Gx����_^[]� �G|�����    �D��6�@�@�Ѓ��    �G|_^[]� �V������W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������U��QW���d �G`t~S�];_xttV�7�ΉE�u��Ǻ���xP u����#��赺���M�S�u�pPj�GP蠺���H ��ЉG|^��u�E�_x��t�    �G`[_��]� �M�Gx������t�3�[_��]� �����������U��E��t	�Ap� �yd t�Ah]� 3��y|��]� ���U���u �D��u�u�@�u�u�@�u�uQ�Ѓ� ]� ���U��D��uQ�@�@�Ѓ�]� ����̡D�Q�@�@��Y�U��D��u�u�@Q�@�Ѓ�]� �̡D��@� ������U��D�V�u�@�6�@�Ѓ��    ^]���������������U��VW���T����u���u�x@�u�A����H ���_^]� ����U��VW���$����u���u�xD�u�����H ���_^]� ����W��������xH u3�_�V�������ύpH�ܸ���H �^_�����U��W���Ÿ���xL u3�_]� V��谸���u���u�pL�u蝸���H ���^_]� U��W��腸���xP u���_]� V���o����u���u�pP�u�u�Y����H ���^_]� ������������U��W���5����xT u���_]� V�������u���u�pT�����H ���^_]� ��U��W��������xX u���_]� V���߷���u�ύpX�ҷ���H ���^_]� �����U���SVW�}�م�t.�M��������蟷���ˍpL�E�P葷���H ��ЍM�� ����u��tW�D��M�Q�@�@�СD��M�VQ�@�@�СD��M�Q�@�@�Ѓ����;����H@��t�D�VQ�@�@�Ѓ�_^[��]� ���������U��VW�������u�΍xH������H ���_^]� ����������U��W���ն���x` u
� }  _]� V��轶���u�ύp`谶���H ���^_]� ���U��SVW��蓶���x` u� }  �#�������ύp`�E���P�l����H ��Ћ��D��]S�I�I�у�;�>�D�S�@�@�Ѓ�;�)���.����u���u�pDS�u�����H ���_^[]� _^�����[]� U��W��������xP u
�����_]� V���ݵ���u���u�pP�u�u�u�u������H ���^_]� ����U��W��襵���xT u
�����_]� V��荵���u���u�pT�}����H ���^_]� U��W���e����xX tV���W����u�ύpX�J����H ���^_]� �������������U����E��E�    P�u�E�    �E�    �E�    �E�    �E�    ��o ����t(�M��t!�u��D��u��u��@�u�Q�@X�Ѓ���]�3���]����������������U��USV��F�����N;�~}��@�+�W�����ρ�  �yI���Au��u	�   +���D�h@�h�   �H��    P�6��  �ЋЃ���t�N�~_�^���^[]� �F_�F��^[]� �^^[]� ��������������U��M�]�`����U��M�]�`����V��h��Vh�����F    �D�h ��@P� �Ѓ��F��^����������̃y ���u�D��q�@P�@��Y���U��I��u3�]� �D�j �u�@P�uQ�@�Ѓ�]� ���U��I��t�D��uQ�@P�@�Ѓ�]� ��������������U��I��t�D��uQ�@P�@�Ѓ�]� ���������������    ���A    �V����t&�D�Q�@P�@L�СD��6�@P�@<�Ѓ��    ^����������������U��SVW�����t�D�Q�@P�@<�Ѓ��    �G    �M�]h���O�D�Sh�h ��@PQ�u�@8��3����9u~E���x u�@   �D��HP���p�A�Ѓ��D�V�7�@P�@@�Ћ���F�A;u|�3�9_^��[]� �����������U���u�E�u�p�,���]� ��������U��SVW��3�9w~=�]�D�V�7�@P�@@�ЋЃ���t-�D�j Sj�APR�@�Ѓ���tF;w|�_^�   []� �D��7�@P�@L�Ѓ�3�_^[]� ������������̡D��1�@P�@D�Ѓ��������������̡D��1�@P�@H��Y���������������̡D��1�@P�@L��Y���������������̡D��@P�@P�����U��D��@P�@T]����������������̡D��@P���   ��U��D��@P���   ]��������������U��M�]�`����U��V��~ ���u�D��v�@P�@�Ѓ��Et	V��������^]� �����������A    �A    �A    ���V��~ ���u�D��v�@4� �Ѓ��F    �F    ^���������������̸   ����������̸   �����������3�� ������������ �������������U��D�V��h�  �@4�v�@$���u�D��u�u�@4�u�v�@�Ѓ�2�^]� ���������������U���u��u�u�u�P]� ��������3�� ����������̸   � ��������� �������������U��Q�D�SVW�@�ً}3��ω]��@ ��=INIb�  ��   =SACbmt)=$'  t
=MicM�f  ���W�P$�   _��^[��]� ��MQ�M��u�Q�ˉu�P��t�D��u�u��@4�s�@�Ѓ��   _��^[��]� =ARDb�  �D���j j�@���   �Ћ؋ϡD�j j�@���   �ЋM���D�j j�@���   �ЋM��D�j j�@���   ���u�M�PVW�S�R�   _��^[��]� ����P�   _��^[��]� =NIVb_tF=NPIbt.=ISIbuV�3���  P���r  P���V�   _��^[��]� ���W�P_^[��]� ����P�   _��^[��]� =cnyst_��^[��]� �D���j hIicM�@���   �Ћ��WP�R _^[��]� �������U���,V��~ t~�D��v�@4�@�Ѓ} t�D�P�F�I0�p�Al�Ѓ�^��]� ���E��M��E�    hARDb�����NP�E�P�E�P�1  �D��M�Q���   � �Ѓ��M�����^��]� ������������U��D��u�q�@4�@l�Ѓ��   ]� �������������̡D��q�@4�@�Ѓ�������������̡D��q�@4�@�Ѓ�������������̡D��q�@4�@�Ѓ�������������̡D��q�@4�@|�Ѓ�������������̡D��q�@4���   �Ѓ�����������U��D��u�q�@4�@(�Ѓ�]� ���U���u�D��u�u�@4�q�@,�Ѓ�]� �������������U��D��u�u�@4�q�@0�Ѓ�]� �D��q�@4�@4��Y���������������U��D��u�q�@4���   �Ѓ�]� U��D��u�q�@4�@ �Ѓ�]� ���U��D��u�q�@4�@$�Ѓ�]� ���U��D�V�uW���   ��V�@�Ѓ����D�V���   u �@@�ЋD�P�w�I4�A �Ѓ�_^]� �@�Ѓ����D�u'���   V�@8�ЋD�P�w�I4�A$�Ѓ�_^]� �@h��h
  ��0  �Ѓ�_^]� ����������U��D��u�u�@4�q�@D�Ѓ�]� U��D��u�u�@4�q�@H�Ѓ�]� U��D��u�u�@4�q�@L�Ѓ�]� U��D��u�u�@4�q�@P�Ѓ�]� U��D�SVW���   �ً}W�@�Ѓ����D����   �@��   �uV�Ѓ����D�V���   u6�@@�ЋD���W���   �I@�ыD�VP�s�I4�AP�Ѓ�_^[]� �@�Ѓ����D�u=���   V�@8�ЋD���W���   �I@�ыD�VP�s�I4�AH�Ѓ�_^[]� h��h�  ��   W�Ѓ����D���   ���   �uV�@�Ѓ����D�V���   u6�@@�ЋD���W���   �I8�ыD�VP�s�I4�AL�Ѓ�_^[]� �@�Ѓ����D�u=���   V�@8�ЋD���W���   �I8�ыD�VP�s�I4�AD�Ѓ�_^[]� h��h�  �
h��h�  �@��0  �Ѓ�_^[]� �����U���u�D��u�u�@0�u�q���   �Ѓ�]� �������U��D��u�q�@0���   �Ѓ�]� U��D����E�@0�$�u�u���   �q�Ѓ�]� U���u�D��u�u�@4�u�q�@�Ѓ�]� ����������U���u�D��u�u�@4�u�q�@�Ѓ�]� ����������U���u,�D��u(�u$�@4�u �u�@T�u�u�u�u�u�q�Ѓ�,]�( ��������U���u�D��u�u�@4�u�q��  �Ѓ�]� �������U���u$�D��u �E�u�@4�u����  �D$�E�$�q�Ѓ�$]�  ���������������U��D�h����h����h�����u�@4�uh�����@Th����h����h�����u�q�Ѓ�,]� ����������U��D��u�q�@4�@8�Ѓ�]� ���U��D��u�q�@4�@<�Ѓ�]� ���U��D��u�u�@4�q���   �Ѓ�]� ������������̡D��q�@4�@@�Ѓ�������������̡D��q�@4��  �Ѓ�����������U��D����E�@4�$�q��  �Ѓ�]� ������U���u�D��u�u�@4�u�q�@X�Ѓ�]� ���������̡D��q�@4�@`��Y��������������̡D��q�@4�@d�Ѓ��������������U���u�D��u�u�@4�u�q��   �Ѓ�]� �������U���u�D��u�u�@4�u�u�@\�u�q�Ѓ�]� ����U��D��u�u�@4�q��  �Ѓ�]� �������������U��D��u�u�@4�q�@h�Ѓ�]� U��D��u�u�@4�q��  �Ѓ�]� �������������U��D��u�u�@4�q�@p�Ѓ�]� U���V��M�hYALf�����D�P�v�R4�Bl�Ѓ��M������^��]���������U��QVW�}�M���t�D��Mj j�@���   �Љ�u��t�D��Mj j�@���   �Љ�D��M�VW�@4�q�@p�Ѓ�_^��]� �������U���u�D��u�I�u�@0�q���   �Ѓ�]� �������U���u�D��u�u�@4�u�q�@x�Ѓ�]� ����������U��D��u�q�@4�@t�Ѓ�]� ���U���u�D��u�u�@4�u�u���   �q�Ѓ�]� ����U���u�D��u�u�@4�u�u���   �q�Ѓ�]� ����U����D�S�E�    �ًM�E�    �@W�{j ���   j�ЋM�E��D�j j�@���   �ЉE��M��D�Q�M�Q�@0�w�@`�СD��s�@4�@�ЋD��U�j R�U�I0R�U�R�U�RP�C�p�Ah�Ѓ�,�} _[t(�} t(�M�U�;�~<�E��;�}3�M��U�;�~)�E���} u�M�U�;�~�E��;�}�   ��]� 3���]� ���U���u�E�D����@4�D$�E�$�u���   �q�Ѓ�]� �����U���u�D��u�u�@4�q���   �Ѓ�]� ���������̡D��q�@4���   �Ѓ����������̡D��q�@4��  �Ѓ�����������V��Vh0E���D��@0� �Ѓ��F�F    ��^�����V��N����t�D�Q�@0�@�Ѓ��F    ^������̸   ����������̸   ����������̸   � ��������3�� �����������3���������������� �����������������������������U��D�VW�}��@�ϋ@ ��=NIVb��   ��   =TCAbwtM=$'  t3=MicM��   �D���j hIicM�@���   �Ћ��WP�R_^]� ���W�P_�   ^]� �D���j hdiem�@���   �Ћ��WP�R_^]� =INIbu�~ u�����F   �P_^]� �~ t�����P_^]� =atni@t1=ckhct=ytsdu;����P_�F    3�^]� ����P_^]� �%�  _3�^]� =cnys����_3�^]� ����������U��V��N��u3�^]� �D�j j j �@0j j �u ���   j �ujQ���u�D��u�u�@0�uj �u���   �v�Ѓ�D^]� ����������̋I��u3�áD�Q�@0�@�Ѓ�����̋I��u3�� �D�Q�@0�@�Ѓ�� U���V�q��u�E�p�    ^��]� �E�H��D�Q�u�M��@0RVQ���   �Ћuj PV�    �F    �D����   �I�ыD��E�P���   �	�у�$��^��]� ��������U��D��u�q�@0���   �Ѓ�]� �D��q�@0���   �Ѓ����������̡D�j j j �@0j j j ���   j j j4�q�Ѓ�(�������̡D�j j j �@0j j j ���   j j j;�q�Ѓ�(��������U��D��u�q�@0�@�Ѓ�]� ���U��I��t'�D�j j j �@0j j j �u���   j jQ�Ѓ�(]� �����������U���u�D��u�u�@4�q�@,�Ѓ�]� �������������U��D��u�u�@4�q�@0�Ѓ�]� �D��q�@4�@4��Y���������������U��V�q��u3�^]� �E�H��D�Q�u�@0RV�@�Ѓ�^]� �����������U��V�q��u3�^]� �E�H��D�QRV�@0���   �Ѓ�^]� �����������U��E3�h���h  �P��j ��BRj �u�u�   ]� ���U���$VW���M�htniv������D��M��uhulav�@�@4�СD��M�hgnlfhtmrf�@�@4�СD��M��uhinim�@�@4�СD��M��uhixam�@�@4�СD��M��uhpets�@�@4�СD��M��uhsirt�@�@4�ЋM �u$��  �u�����t,�D�Qh2nim�M܋@�@4�СD��M�Vh2xam�@�@4�ЍE܋�P�u�E�P�S����D�P���   �@8�ЋD����E�P���   �	�у��M�� ���_��^��]�  ������U���$V��M�htlfv�����D��M��E���@�$hulav�@,�СD��M��u,htmrf�@�@4�СD��M��E���@�$hinim�@,�СD��M��E���@�$hixam�@,�СD��M��E$���@�$hpets�@,�СD��M��uDhsirt�@�@4���U0W�f.џ��Dz�E8f.����D{?�D��M܃��@�$h2nim�@,�СD��M��E8���@�$h2xam�@,�СD��M��u@hdauq�@�@4�ЍE܋�P�u�E�P�����D�P���   �@8�ЋD����E�P���   �	�у��M�������^��]�@ ������������U���u,W�j ��$htemf�E$�� �D$�E�D$�E�D$�E�$�u����]�( ���������������U���Mf.���(��%�����D{�Y��^��Uf.8����D{�Y��^��u,W�j ��$hrgdf�E$�� �Y��^��D$�E�L$�T$�$�u�o���]�( �����������U���u,�p�W�j ��$htcpf�E$�� �^��D$�E�^��D$�E�^��D$�E�$�u�����]�( �����������U���0�E�M���u�D��@���   �Ѕ�u��]� SVW��蜔  htlfv�MЋ��}����u���D�fn���ɋy��Y��E��E��$�Κ �]��F�$��� �E�M��]��^E�G,�$hulav�СD��M�hmrffhtmrf�@�@4�Ћu���D�fn���ɋx��Y��E��E��$�Y� �]��F�$�K� �E�M��]��^E�G,�$hinim�Ћu���D�fn���ɋx��Y��E��E��$��� �]��F�$�� �]��E�M��^E�G,�$hixam�СD��M�������@�$hpets�@,�СD��M�j hdauq�@�@4�СD��M�Shspff�@�@4�СD��M��u hsirt�@�@4�ЋM��E�P�u�E�P�����D�P���   �@8�ЋD����E�P���   �	�у��M�����_��^[��]� ������U���$V��M�hCITb�z����D��M��uhCITb�@�@8�СD��M��uhsirt�@�@4�СD��M��uhulav�@�@4�ЍE܋�P�u�E�P�`����D�P���   �@8�ЋD����E�P���   �	�у��M��-�����^��]� ����U��V�q��u3�^]� �E�E�H��D�Q�u �@0���@(�D$�E�$�uRV�Ѓ�$^]� U����E�Vj �u��MP����P�u��������D����E�P�I�I�у���^��]� �����������U��V�q��u3�^]� �E�H��D�Q�MQ�@0RV�@,�ЋM3҃�9U�^]� �������������U��V�q��u3�^]� �E�H��D�Q�u�@0RV�@,�Ѓ�^]� �����������U��V�q��u3�^]� �E�H��D�Q�u�@0RV�@0�Ѓ�^]� �����������U��VW���O����   �E�P�0�D�R�u�@0VQ�@0�Ѓ���tf� t`�E�H��D�Q�p0�E��P�F0R�w�Ѓ���t8���t1�E�H��D�Q�p0�E��P�F0RW�Ѓ���t_�   ^]� _3�^]� ��������������U��QV�q��u	3�^��]� �EW�E�    �H��D�Q�M�Q�@0RV�@8�Ћ�����t:�U���t3�D��uR�A�@�Ћu�����t�D�V�@�@��V�'�������_^��]� ����������U��V�q��u3�^]� �E�H��D�Q�u�@0�uR�@<V�Ѓ�^]� ��������U��E��V���u�D��@���   �Ѕ�u^��]� W���͎  �v����t!�E�H��D�Q�M�Q�@0RV�@0�Ѓ���fnǍM�������Y���D$�E��Y���$�`M _�o �E� ��^��]� �����������U��D����@V��M�Q�@�Ѓ��E���P�u�U�������t�M�E�P�ӕ���D��E�P�I�I�у���^��]� �����U��V�q��u3�^]� �E�H��D�Qj j �@0j j j ���   j Rj1V�Ѓ�(^]� �������������U��D�Vj �u�@��M���   ��h���h  �j j jj P�u���E���^]� U��D�Vj �u�@��M���   ���u$���u j �u�u�uP�u����^]�  �U����D�W�V����M�@�$�u���   ���E8��j �u@�]����D$�E0�$�u,�E$�� �D$�E�D$�E�D$�E��$�u����^��]�< ����U����D�W�V����M�@�$�u���   ��j j ��W��]���$htemf�E$�� �D$�E�D$�E�D$�E��$�u�8���^��]�$ �U����D�W�V����M�@�$�u���   ���Uf.���(��%����]���D{�Y��^��Mf.8����D{�Y��^�j j ��W���$hrgdf�E$�� �Y��^��D$�E��T$�L$�$�u�t���^��]�$ �������������U����D�W�V����M�@�$�u���   ���p�W�j j �����]�$htcpf�E$�� �^��D$�E�^��D$�E�^��D$�E��$�u�����^��]�$ �������������U���0�D�(��V��M�Q�ufE��@�M�Q�M���   ��j �u ���u�o �E��u�E�P�u�u�x���^��]� �U��D���0�@VW���M��@Q�СD��M����@Q�u�MЋ��   Q�M�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�Ѓ��E����uj P�u�����D����E�P�I�I�ыD��A�M�Q�@�Ѓ���_^��]� ���U���dV��M��O����D��MP�u�R�E�P���   ��P�M��ڏ���M�����j j �E�P�M�蒐��P�u�������D����E�P�I�I�у��M��؏���M��Џ����^��]� �������U���P����U�E�V�uW�����t+�D���W��΋@�$R���   ���]��E��E��D��M�W�Q�ufE��M��E��@Q�΋��   �Ћw�o �E��~@f�E؅�u
_3�^��]� �E�E�H��D�Q�u �Mȋ@0���@(�D$�E��$QRV�Ѓ�$_^��]� ���U��V�q3���t)�E�H��D�Q�MQ�@0RV�@,�Ћ���3�9E���D�P�u�Q�M�R0�ҋ�^]� ��������������U��V�q��t!�E�H��D�Q�MQ�@0RV�@,�Ѓ����D��u�u�A�M�@4�Ћ�^]� ������U���V�q��t!�E�H��D�Q�M�Q�@0RV�@0�Ѓ����D����E��A�M�$�u�@,�Ћ�^��]� �������U���(���E�VP�ufE��u������D����E�P�u�Q�M�R@�ҋ�^��]� �����������U���V��W�WfE�~�E�����   �E�H��D�Q�M�Q�@0RW�@0�Ѓ���tx�~��tq�E�H��D�Q�M�Q�@0RW�@0�Ѓ���tN�v��tG�E�H��D�Q�M�Q�@0RV�@0�Ѓ���t$�D��M�Q�u�M�@�@H��_�   ^��]� _3�^��]� ���������U��D����@V��M�Q�@�Ѓ��E���P�u������D����E�P�u�Q�M�R8�ҡD��M�Q�@�@�Ѓ���^��]� ��������������U���,V��M��?����D��M�Q�@�@�Ѓ��E���P�u�m�������u�D��M�Q�@�@�Ѓ�� �E�P�M��Ռ���D��M�Q�@�@�Ѓ��D��M�P�E�P�u�R<�ҍM�貋����^��]� ���������U��� V�qW��E�fE���t%�E�H��D�Q�M�Q�@0�M�QRV�@<�Ѓ����U���t�D��A�M�Q�MR�@H�ЋU���t�D����E��M�@�$R�@,�Ћ�^��]� ���U��E3�Vh���h  ��8�p�   ��RE�3���j ��@Pj V�u�����^]� ��������������U���u �U3��u�:��P�u�u�u�r�u����]� ���U��U3��E4�:��P�u<���D$�E,�$�u(�E �� �D$�E�D$�E�D$�B�$�u�}���]�8 ���������U��E3�W��8�H��Rj ��$htemf�E �� �D$�E�D$�E�D$�$�u����]�  ������U��E3��U�(��%���8�h��f.�����D{�Y��^��Mf.8����D{�Y��^�Rj ��W�$hrgdf�E �� �Y��^��D$�T$�L$�,$�u�v���]�  ��U��E3��p�W��8�P��Rj ��$htcpf�E �� �^��D$�E�^��D$�E�^��D$�$�u����]�  ��U��U3��:��P�u�B�u�uP�u�u�����]� �����U��E3��u�8��RP�u�����]� ��������������U���$V��M�hgnrs�Z����E�M��E��D��E�   Qj�@�M܋��   �СD��M�Q���   � �ЋE�M��E����D��E�   Q�@�M�j���   �СD��M�Q���   � �Ѓ��E܋�P�u�E�P�����D�P���   �@8�ЋD����E�P���   �	�у��M��ݫ����^��]� ����U��W�y��u3�_]� �E�EV�H��D�Q�u �p0���E���D$�E�$P�F(RW�Ѓ�$^_]� ���������̡D�j j j �@0j j j ���   j j j �q�Ѓ�(��������U��I��u3�]� �D��u�u�@4Q��  �Ѓ�]� ��U��I��u3�]� �D��u�u�@4Q�@h�Ѓ�]� �����U��I��u3�]� �D��u�u�@4Q�@p�Ѓ�]� �����U��I��u3�]� �D��u�u�@4Q��  �Ѓ�]� ��U���u�D��u�u�@0�u�q���   �Ѓ�]� �������U��D��P0�E�pj j j �u�uj �0���   j=�q�Ѓ�(]� �����������U��D��P0�E�p�uj j j��uj �0���   j=�q�Ѓ�(]� �����������U��E����u��EСD��2�@0�u�q�@@�Ѓ�]� �U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�u�u���   �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�u�u���   �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   �u�ujQ�ЋE���(��]� ���������������U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �uj*Q�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�uj �u���   j	Q�ЋE���(��]� �U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�uj �u���   j
Q�ЋE���(��]� �U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�u�u���   �uj'Q�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�u�u���   �uj,Q�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �uj:Q�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj j j �u�E�    �u�@0j j j)���   Q�ЋE���(��]� ���U��Q�I��u3���]� �D��U�Rj j �u�E�    �@0j �u���   j j j)Q�ЋE���(��]� ���U��I��u3�]� �D�j j j �u�@0�u�u���   j �ujQ�Ѓ�(]� ��U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �ujQ�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj �u�E�    �u�@0�u�u���   j �uj>Q�ЋE���(��]� U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U��D�j j j �u�@0�u�u���   j �uj.�q�Ѓ�(]� �������������U��V�q��u3�^]� �E�H��D�Qj j �@0j j �u���   �uRjV�Ѓ�(^]� �����������U��V�q��u3�^]� �E�H��D�Qj j �@0j j j ���   j RjV�Ѓ�(^]� �������������U��V�q��u3�^]� �E�H��D�Q�u�@0RV�@\�Ѓ�^]� �����������U���SVW�u�ٍM��zw���EP�E�P�M��w����tj�}�I �M��tI�D�Q���   �@H�ЋS������tN�w�D�j j j �A0j �u����   V�7jR�Ѓ�(��t"�EP�E�P�M��Pw����u�_^�   [��]� _^3�[��]� ���U��Q�I��u3���]� �D��U�Rj j �u�E�    �u�@0�uj �u���   jQ�ЋE���(��]� �U��D�VW�}��@4�w� �ЋE�G    �w�H��D�Q�u�@0WR�v���   �Ѓ��G3Ʌ���_��^]� �������U��I��u3�]� �D�j j j �u�@0�u�u���   j �uj/Q�Ѓ�(]� ��U��U��u3�]� �r�B    �D��u�q�@0���   �Ѓ�]� ���������U��I��u3�]� �D�j j j �@0j j �u���   j j jQ�Ѓ�(]� ����̡D�j j j �@0j j j ���   j j j6�q�Ѓ�(��������U��I��u3�]� �D��u�u�@0�uQ�@D�Ѓ�]� ��U��I��u3�]�  �u$�D��u �u�@0�u�u���   �u�u�uQ�Ѓ�$]�  �I��u3�áD�Q�@0�@X�Ѓ������U��I��u3�]� �D��u�u�@0Q�@L�Ѓ�]� �����U��Q��u3�]� �D��H0�E   �P�APR�Ѓ�]� ��U��I��u3�]� �D��uQ�@0�@P�Ѓ�]� ��������U��I��u3�]� �u�D��u�u�@0�uQ�@T�Ѓ�]� ���������������U���VW���M��Ν���E�M�P�0�D�RQj �@0j j j ���   j Vj8�w�Ћ���(��t�M�E�P������M�����_��^��]� ����������U��EV�P�0�D�R�u�@0j j j ���   j j Vj9�q�Ѓ�(^]� ��������U��EV�P�0�D�R�u�u�@0�u�u�@hV�q�Ѓ�^]� ��������������U��QVW�}�M���t�D��Mj j�@���   �Љ�u��t�D��Mj j�@���   �Љ�D��M�VW�@0�q�@`�Ѓ�_^��]� �������U���u�D��u�u�@0�q���   �Ѓ�]� ����������U��D��U�@0��t*���   R�q�ЋD����uR�A0���   �Ѓ�]� �u�@|�q�Ѓ�]� ��U���u�D��u�u�@0�u�u�@p�q�Ѓ�]� �������U���u�D��u�u�@0�u�u�@d�q�Ѓ�]� �������U��D�j j �u�@0�u�u���   �uj �uj3�q�Ѓ�(]� ������������U��Ej j j ��D�j j j �@0j Rj�q���   �Ѓ�(]� �������������U��Ej j j ��D�j j j�@0j Rj�q���   �Ѓ�(]� �������������U��Ej j j ��D�j j j �@0j Rj�q���   �Ѓ�(]� �������������U��EV�P�0�D�Rj j �@0j j j ���   j Vj"�q�Ѓ�(^]� ���������U��EV�P�0�D�Rj j �@0j j j ���   j Vj5�q�Ѓ�(^]� ���������U��EV�P�0�D�Rj j �@0j j �u���   j Vj<�q�Ѓ�(^]� ��������U��D�Vj j �@0��j j j �u���   j �uj�v�СD��u�v�@0�@t�Ѓ�0^]� �������̡D�j j j �@0j j j ���   j j j�q�Ѓ�(��������U��D�j j j �@0j j j �u���   j j�q�Ѓ�(]� �D�j j j �@0j j j ���   j j j�q�Ѓ�(��������U��D�j j j �@0j j j ���   j �uj�q�Ѓ�(]� U��D�j j j �@0j j j �u���   �uj&�q�Ѓ�(]� ��������������̡D�j j j �@0j j j ���   j j j(�q�Ѓ�(�������̡D�j j j �@0j j j ���   j j j#�q�Ѓ�(��������U��D�j j j �@0j �u�u���   j �uj+�q�Ѓ�(]� �������������̡D�j j j �@0j j j ���   j j j0�q�Ѓ�(��������U��D��u�q�@0���   �Ѓ�]� U���V�u ��M��̗���D��M��uh8kds�@�@4�СD��M Q�M��E     Q�@0j �u�u���   �u�u�uj2�v�Ћu �M��(著����^��]� �������̡D��q�@0���   �Ѓ�����������U��I��u3�]� �D�j j j �@0j j j ���   j �uj-Q�Ѓ�(]� �����U����D�Wj ���M�@j���   �ЋM�E��D�j j�@���   �ЉE��M��D�Q�M�Q�@0�w�@`�СD��U��H0�E�pR�U�R�U�R�U�R�0�Ah�w�Ѓ�(�} _t(�} t(�M��U�;�~<�E��;�}3�M��U�;�~)�E���} u�M��U�;�~�E��;�}�   ��]� 3���]� �����U��SV�uW��u�q�D��]��j hdiuM�@���   �Ћ���tI;>u	_^3�[]� �D���j hIicM�@���   ��;�u�D���j h1icM�@���   �Шu��>_^�   []� ���������U��D���(�@V�u��hfnic�@T�ЋЅ�t�D�j
�A�ʋ��   �Ѕ���   �D��M�hfnicQ�΋@�@P��P�M��.����M��F����u�E�P���H����M��0����D��΋@�@ �Ѓ��t�D��΋@�@ �Ѕ�u�D���hfnic�@�@$�СD����uj
�@�@8��^��]������������̡D��q�@0���   �Ѓ�����������U���$V��M�hmnrs�Z����D��M��uj�@�@4�ЍE܋�P�u�E�P�s����D�P���   �@8�ЋD����E�P���   �	�у��M��@�����^��]� �������U���$�DSSS�} V��SSSSE��M�P�͓���D��M܋@�@ �ЋD�jP�Q�M܋B4�ЍE܋�P�u�E�P������D�P���   �@8�ЋD����E�P���   �	�у��M�褓����^��]� �����������V��Vh0E���D��@0� �Ѓ��F�F    ���4��F   �F    ^�V��N����t�D�Q�@0�@�Ѓ��F    ^�������U��V��N�F    ��tg�D�j j j �@0j j j ���   j j jQ���u�D��u�u�H03�9E�u����
j P�v���   �Ѓ�D��t�~ t
�   ^]� 3�^]� ��������������U��E�A�I��u3�]� �D�Q�@0�@�Ѓ�]� �����U��D�S�]V�@��ˋ@ ��=ckhc��   t|=cksatb=TCAb��   �D���Wj hdiem�@���   �Ћ��SW���F   �R�~ ��t��t��u3��΃���P�J���_^��[]� �~ ti����P^[]� �~ tV�D�j j j �@0j j j ���   j j j �v�Ѓ�(��t*�F    �   ^[]� =atnit�u��S�x���^[]� ^3�[]� ����������U��Q�y �M���   S�]V�uW�}��wp�$�H29u��   �^9u��   �S9u��   �H9u��   �=�E;�~6;���   �,�E;�|%;�~}��E;�|;�|p��E;�~;�~c�9uu\�D�j j j �@0j j j ���   j �uj�q�Ѓ�(fn����j���D$fn�����$S�o�  �E����@    _^[��]� �y1�1�1�1�1�1�1�1�1����U��W��� �6  V�u����   �$��3�Ef/E�  �   �Ef/E��   �   �Mf/M��   �   �Mf/M��   �|�Uf/Uvp�E f/���   �_�Uf/UrS�E f/���   �B�Uf/Ur6�E f/�w�)�Uf/Uv�E f/�sf��Ef.E���DzT�D�j j j �@0j j j ���   j �uj�w���E ��(�u(���D$�E�$V���  ���G    ^_]�$ ��2�2�2�2�23383Q3U���E j���D$�E�D$�E�$�u�u�]���]�  ���������U���E j���D$�E�D$�E�$�u�u����]�  ���������U���E j���D$�E�D$�E�$�u�u�����]�  ���������V��Vh0E���D��@0� �Ѓ��F�F    ���\��F   ^��������V��N����t�D�Q�@0�@�Ѓ��F    ^�������U��D�V��M�@�@ ��=cksat]=ckhct�u���u�o���^]� j j j j j �F   �D�j j j �@0j �v���   �Ѓ�(��t#�F    �   ^]� �~ t����P^]� 3�^]� �������������U��V��Vh0E���D��@0� �ЋM���F�E�F    �F   ����F�D�j hmyal�@���   �ЉF��t��t�F    �D��Mj
hhfed�@���   �ЉF��^]� U��D�V��M�@�@ ��=ytsdt�u���u����^]� �D��v�@0���   �Ћ�����P�   ^]� ����������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U���V�u�V�E�    �    �B    ������D��E�    j ���   �E�PR�I�ыD��E�P���   �	�у���^��]� ����������̋A��uË ���������������������U��V���PD��t�E9Ft
�F�΋�PH^]� ���������̋A�������������U��j0�u�3y  ��]���������������U��j0�u���  ��P�
y  ��]������U����E�j0�u�uP���  ��P��x  �D��M�Q�@�@�Ѓ���]���������U����E�j0�u�u�uP���  ��P�x  �D��M�Q�@�@�Ѓ���]������U��j$�u�sx  3Ƀ�������]�����U��j$�u��  ��P�Jx  3Ƀ�������]������������U����E�Sj$�u�uP��  ��P�x  �D�3ۃ��E�P�ËI�I�у���[��]������������U����E�Sj$�u�u�uP��  ��P�w  �D�3ۃ��E�P�ËI�I�у���[��]���������U��D��u�u�@j ���   �Ѓ�]�U��D��u�u�@�uj ���   �Ѓ�]��������������U��D��@���  ]��������������U��D��@0���   ]��������������U��D��M����@0VW�u���   �uQ�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]��������������U���4�D�SV�u�@WV�@�СD����M3ۋ@SS���   �ЋM�E��D�Sj�@���   �Ћ����M  3ɉM�d$ ��~k�D��M�Q�@�@�СD��M�j j�h��@Q�@�СD����΋@�@<�ЋȍU�D�j�j�R�@Q�΋@L�СD��M�Q�@�@�Ѓ��D��M�W�u��@0Q���   �Ћ��MܡD�Q�@�@�СD��M�QW�@�@�СD��M�Q�@�@�СD����΋@�@<�ЋȍUܡD�j�j�R�@Q�΋@L�СD��M�Q�@�@�СD����MC��
�M�@j Q�M���   �ЋM�E�A�D�j Q�M�P���   �ҋ��������_��^[��]����U��D��@0���   ]��������������U��D��@0���   ]��������������U��D��@0���   ]�������������̋�W�R�J��A(�P$j j h����x  �������������̸������������U���(V��M�WQ�΋�P(�V����t&�D�j j j �A0j j j ���   Wj jR�Ѓ�(�D��M�Q�@�@�СD��M�Q�@�@�ЋN����t&�D��U�j j j �@0Rj j���   j?j Q�Ѓ�$�D��M�Q�@�@�СD��M�Q�@�@�ЋN����u3��:�D��U�Rj j j h  
 j�U��E�    �@0Rh�  j���   Q�Ћ}���(�D��M�Q�@�@�Ѓ���u_3�^��]áD��M�Q�@�@�ЋN����t&�D��U�j j j �@0Rj j ���   j8j Q�Ѓ�$�D��M�Q�@�@�ЋN����t�D�jQ�@0�@P�Ѓ��D��M�Q�@�@�Ѓ��M�赃��Ph   h  K j;�E��Ph	��h�  ������D��M�Q�@�@�Ѓ��M��׃���N��t�D�Q�@0�@X�Ѓ��N��t�D�Q�@0�@X�Ѓ��N��t&�D�j j j �@0j j j���   j j jQ�Ѓ�(j�v$�pq  ���   _^��]���U���V��Wj�N�\����F4    W��F8    �F<    �F(�D�h�   �v�@0�@�СD��M�Q�@�@�СD��M�j j�h,��@Q�@�Ѓ��E��  �E��E�    ��j j P�E�P������D��M�Q�@�@�Ѓ��Nj j若��_^��]������U���\�D�VW���Mȋ@Q�@�СD��M�j j�h0��@Q�@���G(�Yp��D��E��  �E�    �@�,ȋ@(Q�M�Q�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M��8�@�@<�ЋD�j�j��Q�M�QP�M�BL��j j �E��P�E�P������D��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ��M�htats�����D��M�jj�@�@0�СD��M��G(���@�$j�@,�ЍE��E��  P�E��E�    P�E���P�����D��M�Q���   � �Ѓ��4 t_�D��O0�@P�@h�ЋG4��t�w8�Ѓ��G<�G8    �G4    ��D�h��h�  �@��0  �Ѓ��D��O0�@P�@l�ЍM�肀��_^��]� ����������U��D���@�@VW�}��@ ����=MicMtc=ckhctG=fnic��   j�M������MP�8����M�� ����D��Mjj�@�@4��_�   ^��]� ����P��_���^��]� �D���j hIicM�@���   ��=���uhtats�M��}���D��M�j j�@�@0�ЍE��E��  P�E��E�    P�E��P舸���D��M�Q���   � �Ѓ��M��j���N�F   ��t�D�Q�@0�@�Ѓ��u��W�����_^��]� ��������U��mV��t3�^]� j�N�#���j�m  �N���F    ��t�D�Q�@0�@�Ѓ��   ^]� j������j��l  ��3�����������U���E�A(]� ��������������̍A�������������U��VW��~4 t@�I �D�h��h~  �@��0  ��j
�Ox  �D��v �@P�@�Ѓ���uM9F4uáD��N0�@P�@h�Ѓ~4 t:�D�h��h�  �@��0  �СD��N0���@P�@l���r���_3�^]� �E�N0�F8�E�F4�D�S�@P�@l�Ѓ~4 t#j
�w  �D��v �@P�@�Ѓ���u99F4uݡD��N0�@P�@h�Ћ~<�N0�F<    �D��RP�Rl��[��_^]� [_3�^]� U����M�V�}���M�D���t �@4Q�@�Ѓ���t$��M�Q�u���R(�1�@0�u�@�Ћȃ���u�M�3��}����^��]Ë�U�R�u�P ���M�D��@�@ �Ѓ��t�D��H0�E�P�u�Ix�у��M���|����^��]��������U��D�Vj �u�@��M���   �Ћ���u�    �F^]� ��u9Ft�   ^]� ���������U��V�uW��;uuz�D��Mj htsem�@���   �Ѕ�u\�D��Mj hrdem�@���   �Ѕ�u>�E�E�H��t1�D��Uj RV�@0Q�@,�Ѓ���t�u���  _�   ^]� _3�^]� ���������������U��D���@�@VW���M��@Q�СD��M�Q�@�@�СD��MЃ��@Q�u�M����   Q�M�ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�СD�����@V�@�СD��M�VQ�@�@�Ѓ����%  �D��M�Q�@�@�Ѓ�_^��]� ���������U���SV�u��;u��   �D��Mj htsem�@���   �Ѕ���   �D��Mj hrdem�@���   �Ѕ���   �D��M�Q�@�@�ЋM�E���u��E�    P�E�P�8�����u3��4�D�����@V�@�СD��M�VQ�@�@�Ѓ����A  �   �D��E�P�I�I�у���^[��]� ^3�[��]� ���U��D�Vj �u�@��M���   �Ћ���u�    �F^]� ��u9Ft�   ^]� ���������U���V�uW��;uup�D��Mj htsem�@���   �Ѕ�uR�D��Mj hrdem�@���   �Ѕ�u4�M�E�E��EP�E��u�P虼����t�u���  _�   ^��]� _3�^��]� ����U����D�W�V����M�@�$�u���   �Ћ�]����u�E��    �F^��]� ��u�Ff.E����D{�   ^��]� ����U���SV�u��;u��   �D��Mj htsem�@���   �Ѕ�um�D��Mj hrdem�@���   �Ѕ�uO�EW��E��H��t=�D��U�j RV�@0Q�@0�Ѓ���t!�E������$�,  ^�   [��]� ^3�[��]� �����U���H�D�W�V���E��M�Q�ufE�@�M�Q�M���   ���o �~H��EЃ��u�F�    f�N^��]� ��u5�Ff.EП��Dz�Ff.E؟��Dz�Ff.����D{�   ^��]� U���4�ES�]�M�V�uW�};�t;�t;���   �D��Mj htsem�@���   �Ѕ���   �D��Mj hrdem�@���   �Ѕ�ui�MW��E��E��E�E�P�E��E�P�E�u�P�E�}�PfẺ]�������t.�oE̋M������ �~E�f�@��  �   _^[��]� _^3�[��]� ����U��� �D�(��V��M�Q�ufE��@�M�Q�M���   ���o ��E����u�    �F^��]� ��u�E�P�FP��   ����t�   ^��]� ������U���SV�u��;u��   �D��Mj htsem�@���   �Ѕ�ui�D��Mj hrdem�@���   �Ѕ�uK(���M�E��E�P�u�E��u�PfE��)�����t"�oE���ˋ�� �0  �   ^[��]� ^3�[��]� ���������U���V�uW�}�f.���Dz�Ff.G���D{Y�G���Y��E��E��$�P �F�Y�]��E��E��$��O �E����]�f.E����D{_�   ^��]�_3�^��]����U��V��~ ���u�D��v�@4� �Ѓ��E�F    �F    t	V��L������^]� ��������U��V��N����t�D�Q�@0�@�Ѓ��E�F    t	V�L������^]� ���������������U�����u�E�    �A]� ��u�A;Et�   ]� U�����u�E�    �A]� ��u�Af.E���D{�   ]� ����U�����u�oE�    �A�~Ef�A]� ��u6�Af.E���Dz �Af.E���Dz�Af.E���D{�   ]� ����������U��V�����u�oE�    �F^]� ��u�EP�FP��������t�   ^]� �����������U��V�����u �    �D��P�FP�EP�B�Ѓ��"��u�D��MQ�N�@�@x�Ѕ�t�   �D��MQ�@�@�Ѓ�^]� ��������U��D��@ �@h]�����������������U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��D��uQ�@ �@�Ѓ�]� �����U��D��uQ�@ �@�Ѓ�]� ����̡D�Q�@ �@��Y�U��VW�}����?q���D�WV�J �I�у���_^]� ����U��D��uQ�@ �@ �Ѓ�]� ����̡D�Q�@ �@,�Ѓ���������������̡D�Q�@ �@0�Ѓ����������������U��D��uQ�@ �@4�Ѓ�]� ����̡D��@ � ������U��V�u���t�D�Q�@ �@�Ѓ��    ^]��������������������������U��D���� V��W�}��~D�F<    �F8    �F@    �FH    �FL   �FP    �FT    ����   �E��P�#B  P�N�O���M���K�����E  �F�ύE�P�]M  W�o �F�D��@@�@,�Ћ�����tH�D�j h6  �Q�ϋ��   �҉FP�ϡD�j h5  �@���   ��_�FT^��]� �F   _^��]� ������������̋I@��t�D�Q�@�@D�Ѓ�ø   �̡D��@���   ��U��D�V�u�@�6���   �Ѓ��    ^]�����������̡D�Q�@���   ��Y��������������U��EWɋMW�HH H0H@HP� (���@(��f�H�@0f�H(W�f�H@����@Hf�HX�o� �~Af�@]�������U��EWɋMW�HH H0H@HP� (���@(���@0f�H(W�f�H@f�H����@Hf�HX��@�A�@8�A�@X]������������U���W�W�V�uNN N0N@NP�(���F(���F0W�f�Nf�N(f�N@����FH�Ef�NX��4 �E��E��D �U�f(�fW`����VX�N@�FP�V8^��]�����U���W�W�V�uNN N0N@NP�(���F(���F0W�f�Nf�N(f�N@����FH�Ef�NX�O4 �E��E�@D �U�f(�fW`����V�NH�F(�VX^��]�����U���W�W�V�uNN N0N@NP�(���F(���F0W�f�Nf�N(f�N@����FH�Ef�NX�3 �E��E�C �M����F0fW`��N�F �N8^��]���������U������   V�u�V �F(��^(�Y��Y��X�(��Y��X���D f(�W�f.џ��Dz2W�fD$X(��D$P�D$h�D$`�D$8�D$X�D$�K����^��N�Y��L$�L$X�N �Y��L$8�L$`�N(�Y��L$P�L$h�N0�^8(��V@�Y�(��Y��X�(��Y��X��3D f(�W�f.џ��Dz#W��L$0f�$�   ��$�   �D$@�E����^��N0�Y��L$@��$�   �N8�Y���$�   �N@�Y��L$0�fP�VH(��^X(��Y��Y��X�(��Y��X��C f(�W�f.џ��Dz$W��L$fD$x��$�   f(��L$x�<����^��NH�^P�VX�Y��Y��Y��L$x��$�   �T$�E��$�   �\$p�L$H����  �$�T`�D$0��fW`��$��/  ���\$�D$��0 fW`�fTP�f/�v6�D$h݄$�   �cW �\$ ݄$�   ݄$�   �LW �\$(�D$(��  �D$`W��D$X�D$�'W �D$0f/���\$ ��  �@��\D$ �D$ �  �D$@���$�9/  ���\$(�D$(�D$�10 fTP�f/�vR�D$0fW`��D$�D$݄$�   �V �T$HfW`��\$�T$�D$�D$X�pV �\$ �  �D$hW��D$�D$8fW`��D$�D$�=V W�f/D$@�\$ ��  �(��\D$ �D$ �  ��(�fW`��$�O.  ���\$ �D$ �M/ fTP�f/�v6݄$�   �D$X��U �\$(݄$�   ݄$�   �U �D$(�\$�C  W��D$�D$8fW`��D$�D$݄$�   �rU W�f/D$H�\$�	  �D$fW`��D$��  �D$8��fW`��$�-  ���\$(�D$(�D$�y. fW`�fTP�f/�v-�D$h�D$X��T �\$ ݄$�   ݄$�   ��T �\$�v  �D$xW�݄$�   �D$ �T �D$8f/���\$�E  �D$�X(��D$�,  �D$P���$��,  ���\$ �D$ ��- fTP�f/�vB�D$8fW`��D$�D$�D$X�*T �D$0fW`��\$(�D$�D$�O����T$HW�fW`�݄$�   �T$�D$�D$��S W�f/D$P�\$�s  �D$�\(��D$�Z  ���$��+  ���\$�D$��, fTP�f/�vE�T$HfW`��T$�D$݄$�   �[S �D$8fW`��\$ �D$�D$�����݄$�   W��D$X�D$�!S W�f/D$p�\$ ��  �D$ fW`��D$ �  (��Y�f(��Y��X��> �h�f(�f/��l$@��   �T$8W��\$P�Y�f(��Y��L$�XT$�X�f/��r�L$�5���f/�r�(��D$�(��# �\$PW��D$�d$pf/�v���f/�����f/��D$ ��  �@��\D$�D$�  �\$W�f/��(��T$H�L$�^�v^f/��r���fW`��   ���f/�r���fW`��l(��Q �l$@f(�fW`�W��Mf/��r
����5���f/�r
����(��aQ �(�f(��l$@W��X�f/��T$�T$0v�X@��T$0�T$�d$p�^�(��P' �D$ �D$0�O* �D$@�D$0�>: �\$@W��L$8�Y\$�YD$P�Y��X��X�f/��rf(��#���f/�r
�(��(��! W��D$�L$8f/�v�@��\�f(��D$�E�oD$^�L$� f�H��]ÍI �X�YyZ�\D[\����U������V�uW�W�}��W�F(��Y�(��Y��X��; �h�f(�f/��T$v<�GW�f/���v(���f�N_^��]�(���f�N_^��]��Gf/����^�vTf/��r���fW`��z���f/�r���fW`��Z(��EO �T$fW`��Bf/��r
����&���f/�r
����(��O �T$�X(���G�^��!% �F��W�_�F^��]�������������U���   V�uW��f.��E���D��   �Ff.����Dzq�Ff.����Dzb�EW�^HH H0H@HP� (���@(���@0f�HW�f�H(f�H@����@Hf�HX��]��E�W�}�[7 ��u7�E���H' �E��F�97 f(��F�M��&' �E��5f(���M��' �E��F��6 �E��F��& �E��F��6 �E��F��& f(���p������  �$�`h�m�E��e�f(��YU�f(�P�}�f(��YǍE�Pf(��YߍE��Y��Y��\�f(��Y��M�f(��X��Y��Y��U��U�f(��YE��E�f(��Ye��Y��\��E�f(��Y��Y��]��E�f(��YE��U��X��M��  �m�f(��YE�f(��YU�f(��}�fW`��E�f(��YE�f(��YM��Ye��Y��X��m��E��YE��M�(��YM��\��U��E�f(��Y��E�f(��Y�fW`��E�f(��Y��YU��Y��X��   �e�f(��E�f(��m��M��}��Y��Y�fW`��E�f(��Y��E�f(��Y��E�f(��Y�f(��Y��Y��E�f(��Y��X�f(��Y��M�f(��\��Y�f(��Y��Y��U��Y��X��Yu��E�P�\��eЍE�P�u��E��M��  �e؍E��m�f(��}�f(��Y�f(�P�YE��E�P�YߍE�f(�fW%`��YM��YU��e��\�f(��Y��M�f(��YM��E�f(��YE��X�f(��Ym��U��U��Y��Y��X�f(��Y��\��M��E�f(��YE��Y��]��E��u���   �}��E��e�f(��YU�f(�P�m�E��Y�f(�P�Y]��E�f(��Y��Y��\�f(��Y��M�f(��X��Y�(��Y��U��U��Y��Y��E�(��Y��Y��X�f(��Y�fW%`��Y��\��M��e��u��E��E��E�fW-`��m��MW�P��x����]�W�Pf�x����$!  �E_^��]��e�f(��YM�(ċE�YE�f(�_�m���p���f(��YM�f(�^fW`��Yu��Y]��E��YU�f(��YE��Ym��Y}��X���p���(��\�f(��Ye��YM�f(��YE��Y]�f��\��E��YE��X�W�fW`�XX X0X@XP�E�W�� �E�f��oE��H�M�f��p0�@Hf�Xf�P(f�h@f�xX��]Ë�;c�c�dEg|eLf��������U�������   V�uW�o�o^ �oV��$�   �oF0f���$�   �oF@f(���$�   �oFP�Y���$�   f(��Y��T$ (�f��X�f(�)T$P�Y��X��2 W�f.����Dz)W��L$PfD$ �D$(�D$�D$ �D$8�7����^�f(��YD$ �D$8f(��YF �YL$P�D$�L$P��$�   ��$�   (��Y���$�   �Y��X�(��Y��X��2 W�f.����Dz,W�fD$ (��D$�D$(�D$@�D$ �D$ �A����^�f(��Y�$�   �D$ f(��Y�$�   �Y�$�   �D$@�L$��$�   ��$�   (��Y���$�   �Y��X�(��Y��X��X1 f(�W�f.ʟ��Dz)W�f(�fD$h�D$p�d$h�D$H����9���f(��^�f(�f(��Y�$�   �Y�$�   �Y�$�   �l$H�L$@�XL$8�d$�X��\��Y��f/�s$���f/�r
�(��(�� f(��L$�\L$H�\$�\\$P�u�}f(��L$�Y���T$�\T$ �(��Y��\$�^�T$�X��V(��Y��X��(0 W�f.����Dz	W�f(��<����^��D$�d$�Y��Y��D$h�D$�d$p�Y�fT$h�f�F�f.����Dz2�Ff.����Dz#�Ff.����Dz(���f�N�_^��]��������U���������@W�W�V�uW�}NN N0N@NP�(���F(���F0W�f�N�FHf�N(f�N@f�VX�f.����Dz"�Gf.����Dz�Gf.����D��  �Ef.����D��  �Y���E��, �D$�E�� ��_�D$�G�Y��Y��\$�X�f(��Y��X��v. f(�W�f.˟��DzW�fD$0�|$8�t$0�'����^��7��\$�Y��Y��Y��D$�l$�Y��Y��Y���f(��Y�f(��Y��\$�Y�f(��Y��|$f(��Y��D$(f(��Y�f(��Y��D$(��Y�f(��Y�(��Y�(�����D$ �D$�Y��Y|$�L$0�XL$�D$�X��Xt$ �\�(��\��X�f�����Vf�N(�L$�XL$ �\�(��\L$(�X|$(f��oD$0�n0�\D$f�N@����\�f��FHf�NX_��^��]���������U���p�EV�uW�o�E���wB�$��r�(���F�X��X��\V�=�(��Ff(��\�X���(��f(��\F�X��V�XӋ}���]�f��M��\�U��^@��]��E��$�]��F. �M؃��@��]��\M��Y�f/(�f(��M��X�U�r�\��\��M��U��M����\O�^��M��E��$�M���- �M����@��]��\M��Y�f/(�f(��M��XW�U�r�\��\��M��U��W���~N�\��^��M��E��$�M��a- �MЃ��@��]��\M��Y�f/(�f(��M��XW�U�r�\��\��M��U��]����\�^��]��E��$�]���, �M���@��]��\M��Y�f/(�f(��M��X�U�r�\��\��M��U��U����\W�^��U��E��$�U��, �E����@��]��\E��Y�f/(�f(��E��XW�U�r�\��\��E��U��E����\G�^��E��E��$�E��, �M����@��]��\M��Y�f/(�f(��Xg_^r�\��\��P��]�fT��U�fT؋EfT��X��]�fT��X��M�fT��X��]�fT��X�f/�v�oE�� f�`��]��oE�� �E�f�@��]�#oo>o#oo>o����U����M�Q�	(��Y�Y��Y��X�(��Y��X�W�f.��M����Dz�E �@��]ËU�E�B�p�8�\���j�\��`f(��\̋E�Y���Y��Y�X�(��Y��I�X���^U��Y��Y��Y��X���X��X��\��\�� �B�\��h�@��]�������������U��E�M�p�f(��yf(��!�X�i�Y̋E�Y��X�f(��Y��X��Y��Y��Y��Y��\��\��\�� �x�h]���������U�������   ��3ĉ�$�   �MW�SVW�}�o��oA�G�oA �G �oA0�G0�oA@�G@�oAP�GP�Gf.����Dz%�G f.����Dz�G(f.����Dz�   �3��G0f.���$�   ���Dz%�G8f.����Dz�G@f.����Dz�   �3��GHf.���$�   ���Dz%�GPf.����Dz�GXf.����Dz�   �3���$�   ��H��   H��   H��  (��W�(���D$HW�f�L$@�D$x�oD$@��Gf�L$X�oD$Pf�L$p����G �oD$p�W0f֌$�   �G@�o�$�   �m  3��I ����    t@��|��X  @�����$�@��P�D$<P�>�������  ���  ����   �PW��GXf(��YG8�YW@�_0�gH�\�f(��YG@�Yg8�T$ f(��Y��YWX�\��\��oD$ f��Gf�g(�Gf.����Dz+�G f.����Dz�G(f.����Dz����G����   �(�G �YGX�YP�W�wHf(��YOX�YWP�\�f(��Yw �YG(�\��\�f�W��0f�w@�G0f.����Dz+�G8f.����Dz�G@f.����Dz����G8��$�    ��   �@�G8�YG(�Y �W0�wf(��YO(�YW �\�f(��Yw8�YG@�\��\�f�W��Hf�wX�GHf.����Dz+�GPf.����Dz�GXf.����Dz����GX��$�   ��P�0  �o �M��o@�G�o@ �G �o@0�G0�o@@�G@�o@P�GP�   ��$�   �   �D$�T$�; u\���4@�D����T��Y��Y��Y��X��X��5# ��D$�T$f(��D�f�fY��Y���D��M@���D$J�T$u����o ��~@f�G��$�   ��_^[3��� ��]��������������A    ���d   �U��E�A    �]� �������������U����@i�� %����fn�������X����^���E��E���]���U����@i�� %����fn�������X����^���Y��\���E��E���]���U������V��~ �  �-��W��5��%���@i�� ���������fn�����X����Ai�� �^�%����fn�������Y��X����\��^��T$�Y��\�f(��D$�Y�(��Y��X�f/��L$�p���f.˟��D�b���f(��X; �Y���^D$�! f(��F   �YD$�YL$�Yx��N�X���D$�D$^��]��F�x��F    ^�����]����������������U������V��~ �  �-��W��5��%���@i�� ���������fn�����X����Ai�� �^�%����fn�������Y��X����\��^��T$�Y��\�f(��D$�Y�(��Y��X�f/��L$�p���f.˟��D�b���f(��: �Y���^D$�� f(��F   �YD$�YL$�YP��N�D$�D$^��]��F�P��F    ^��]��������������U��E��Hf(�f/��pvf(�f/�vf(�f/�f(�vf(�f/�vf(�W�f/���   f(��=���^��\��p�f/�v�E�h ]�f.�f(��\ş��Dz
�\��^��2f.˟��Dz(��\��^��X���\��^��X0�(��^��f/�v�X���E��x�X]ËE�` ]�������������U���p���V�uf/F��Vv(�(���   f.�����DzW��Y�����M��E��$�M��"  �m����~�%���]��M�f(��\��V�,�f(�f(��Y��\�H�Y��\�f(��\��Y��Y��\��Y��w>�$��~f(�f(��4f(�f(�(��+f(�f(��!(�f(��(�f(�f(��(�f(�f(ӋE^��@�P��]ÍI )~3~@~J~S~��������U��E���(�`f/��pvf(��f(�f/�vf(�f/�vf(��f(�f/�wf(�f(�W��X�f(��Y=��f/��}�r	f(��  f(��\�f/��}��}�r�E�H��]��=��f/}�s���\��\��}�f.ٟ��D{(��^��M�f(�f(��\�f.��^�f(��\��\���^M��^}���Dz"f.����Dz
�X8��d����\��Vf.���Dz)f.���Dzf(��X���4� ��\�(��#f.���Dz(��X ���8��\��^���E��}�E��@�x��]�����������U��E����=���Pf/���`�Y�rf(��X���Y��f(�(��X��Y��\�W�f(��Y-�f.��\���D��  f.�����D��  (��X%��f/�v�\��
f/�v�X����f/��5��vf(��\��Y��^��X��C���f/�vf(��/f/�v%(�f(��\��\��Y�����^��X��f(�f/�(�v�\��W�f/�v(��X�f/�vf(��\��Y��^��X��P�%��f/�vf(��<�%��f/�v*���f(��\��\��Y�����^��X��f(��\��f/�v�\��W�f/�v�X�f/�v#�\͋E��Y��`�^��X��H]��5��f/�wS�5��f/�v'�\͋E�\���`�Y��^��X��H]ËEf(���`�H]�f(�(�E��`�H]�̡D��@���   ��U��D�V�u�@�6���   �Ѓ��    ^]������������U��D�j �u�@���  �Ѓ�]����U��D�V�u�@�6���  �Ѓ��    ^]������������U��D��@���   ]��������������U��D�V�u�@�6���   �Ѓ��    ^]������������U��� �D�W�j j j fE��E�    �E��E�    �H�E�Pj �E�P�EPPP�u��d  �u�u�uj �Ѓ�8��]�����U��D��uQ�@���   �Ѓ�]� ��U���u�D��u�u�@�u�u���   �uQ�Ѓ�]� ���U���u�D��u�u�@�u�u���   �uQ�Ѓ�]� ���U���u�D��u�u�@�uQ���   �Ѓ�]� ���������U���u�D��u�u�@�uQ��  �Ѓ�]� ���������U��D��u�u�@Q���   �Ѓ�]� ���������������U��VW�}����/=���D�WV�J���   �у���_^]� �U��D��uQ�@���   �Ѓ�]� ��U��D��uQ�@��  �Ѓ�]� �̡D�Q�@��0  �Ѓ�������������U��D��u�u�@Q��t  �Ѓ�]� ���������������U���u�D��u�u�@�uQ���  �Ѓ�]� ���������U��U��tA���    t8�MV��  ;q}(��t	�E�    �	��  �t	�E�    ^]�����    ����������V����t�D�Q�@��<  �Ѓ��    ^������������U��V����t�D�Q�@��<  �Ѓ��    �D��u�u�@�u��8  ��3ɉ��������^]� ��������������V����t�D�Q�@��<  �Ѓ��    ^������������U��	��t�D��u�u�@Q���  �Ѓ�]� ���������U��	��t�D��u�u�@Q���  �Ѓ�]� ���������U��D��@��P  ]��������������U��D��@��T  ]��������������U��D��@��X  ]��������������U���V�u����\E�^@��E��E��$�E��� �M����@��]��\M��Y�f/(�f(��M��XE�r�\��\��M���E�^��]�������������U��EW�AA A0A@AP�o ��~@�Ef�A�o �A�~@�Ef�A(�o �A0�~@�Ef�A@�o �AH�~@��f�AX]� ������U���Mf/��r���]����f/�r���]�(��' �E�E]���������������U���@�i �a(f(��y@f(��YA8�E�Y�q0�Y��\�f(��Y��U�f(��Y��\�f(��Y��U�f(��YQ8�\��AP(��E��Y��U��QX(��Y��\�(��Y��M��IH�E�(��Y��e��\��e�(��Y��m�(��Y�(��YY8�Y��\�(��Y��Y��e��\�(��YI8�Y��\�W��\�W�PP P0P@PP��oM�f��E�f����H0�Xf�@@�E�f�Pf�h(�oM�f��E��HHf�@X��]� �������U������V���N�V f(��^(�Y��L$(��Y��T$�\$�X�(��Y��X��� f(�W�f.ȟ��D{9����^��L$�Y��N�L$�Y��N �L$�Y��N(�N0�V8(��^@�Y��L$(��Y��T$�\$�X�(��Y��X��3 W�f.����D{9����^��D$�Y��F0�D$�Y��F8�D$�Y��F@�NH�VPf(��^X�Y��L$(��Y��T$�\$�X�(��Y��X�� f(�W�f.ȟ��D{9����^��L$�Y��NH�L$�Y��NP�L$�Y��NX^��]����������̡D�Q�@L���   �Ѓ�������������U��D��u�u�@LQ���   �Ѓ�]� ���������������U��D�V��V�@L���   �Ћȃ��D���u�@LQ�u���   V�Ѓ�^]� ���   �@P�ЋD�P���   �M�BH��^]� �������������̡D�Q�@L��(  �Ѓ�������������U��D��u�u�@LQ��,  �Ѓ�]� ��������������̡D��@L� ������U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D��@L���   ��U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��D����u�@LQ�M�Q�@�ЋM��P�Y4���M��q4���E��]� ��������U��D��u�u�@LQ�@�Ѓ�]� ��U��D��uQ�@L���   �Ѓ�]� �̡D�Q�@L�@�Ѓ���������������̡D�Q�@L�@�Ѓ���������������̡D�Q�@L�@�Ѓ����������������U��D��u�u�@L�uQ�@ �Ѓ�]� ���������������U��D��uQ�@L��4  �Ѓ�]� ��U��D��u�u�@L�uQ�@$�Ѓ�]� ���������������U���u�D��u�u�@L�uQ�@(�Ѓ�]� �����������̡D�Q�@L�@,�Ѓ���������������̡D�Q�@L�@0�Ѓ���������������̡D�Q�@L�@4�Ѓ���������������̡D�j Q�@L�@8�Ѓ��������������U��D��u�u�@LQ��  �Ѓ�]� ���������������U��D��@L���   ]��������������U��D��@L���   ]��������������U��D��@L��l  ]��������������U��D��@L���   ]��������������U��D��@L���   ]��������������U��D��@L���   ]��������������U��D��@L���   ]��������������U��D��@L���   ]��������������U��D��@L���   ]��������������U��D��uQ�@L�@<�Ѓ�]� �����U��D��@L���   ]�������������̡D�Q�@L�@��Y�U��D��u�u�@LQ�@@�Ѓ�]� ��U��D�j �u�@LQ�@D�Ѓ�]� ���U��D�j�u�@LQ�@D�Ѓ�]� ���U��D�j �u�@LQ�@H�Ѓ�]� ���U��D�j�u�@LQ�@H�Ѓ�]� ��̡D�Q�@L���   �Ѓ�������������U��D����u�@LQ�M�Q��  �ЋM��P��/���M���/���E��]� �����U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �G�  j �E܋�P�E�P�2�����M���蹊  ��t3���D��M�Q���   �@8�Ѓ����D��E�P���   �	�у���^[��]����������U���$V�E��E�   ���E�   P�M��E��  �E�    �E�    計  j�E܋�P�E�P�1���M���  �D��M�Q���   � �Ѓ�^��]�����U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �7�  j �E܋�P�E�P��0�����M���詉  ��t
�M�-	��� �D��M�Q���   �@L�ЋM��P�	���D��E�P���   �	�ыE��^[��]� ���������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    臇  j �E܋�P�E�P�F0�����M������  ��t
�M�}��� �D��M�Q���   �@L�ЋM��P�	���D��E�P���   �	�ыE��^[��]� ���������U���$�D��E�    �E�    V���   ���u�M�Q�@(�Ѓ��E��  �E��E�    �M��E�    P辆  j�E܋�P�E�P�/���M��5�  �D��M�Q���   � �Ѓ�^��]� ��������U���$�D��E�    �E�    V���   ���u�M�Q�@(�Ѓ��E��  �E��E�    �M��E�    P�.�  j�E܋�P�E�P�/���M�襇  �D��M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    跅  j �E܋�P�E�P�v.�����M����)�  ^��[tW��E��E���D��M�Q���   �@<�Ѓ��D��M�Q�]����   � ���E�����]����������������U����E�E�V���E�   P�M�E��E��  �E�    �E�    ��  j�E��P�EP��-���M�|�  �D��M�Q���   � �Ѓ�^��]� ���������������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    臄  j �E܋�P�E�P�F-�����M������  ��t3���D��M�Q���   �@8�Ѓ����D��E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    ��  j�E܋�P�E�P��,���M��`�  �D��M�Q���   � �Ѓ�^��]� ���U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �w�  j �E܋�P�E�P�6,�����M�����  ��t8�D��E܋uW�P���   �����F�	�у���^[��]� �D��M�Q���   �@P�ЋD��u�o ���   �E�P��	�у���^[��]� �������������U���$�D��E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�~�  j�E܋�P�E�P�]+���M����  �D��M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ��  j �E܋�P�E�P��*�����M����y�  ��t8�D��E܋uW�P���   �����F�	�у���^[��]� �D��M�Q���   �@P�ЋD��u�o ���   �E�P��	�у���^[��]� �������������U���$�D��E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P��  j�E܋�P�E�P��)���M�腂  �D��M�Q���   � �Ѓ�^��]� ��������U��D����@Lj�u���   Q�M�Q�Ѓ��o �E� ��]� ������������U��D����@Lj �u���   Q�M�Q�Ѓ��o �E� ��]� ������������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    ��  j �E܋�P�E�P��(�����M���艁  ��t8�D��E܋uW�P���   �����F�	�у���^[��]� �D��M�Q���   �@P�ЋD��u�o ���   �E�P��	�у���^[��]� �������������U���$�D��E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�  j�E܋�P�E�P��'���M�蕀  �D��M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �~  j �E܋�P�E�P�f'�����M�����  ��t8�D��E܋uW�P���   �����F�	�у���^[��]� �D��M�Q���   �@P�ЋD��u�o ���   �E�P��	�у���^[��]� �������������U���$�D��E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�}  j�E܋�P�E�P�&���M��%  �D��M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �7}  j �E܋�P�E�P��%�����M����~  ��t3���D��M�Q���   �@8�Ѓ����D��E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    �|  j�E܋�P�E�P�x%���M��~  �D��M�Q���   � �Ѓ�^��]� ���U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �'|  j �E܋�P�E�P��$�����M����}  ��t8�D��E܋uW�P���   �����F�	�у���^[��]� �D��M�Q���   �@P�ЋD��u�o ���   �E�P��	�у���^[��]� �������������U���$�D��E�    �E�    V���   ���u�M�Q�@,�Ѓ��E��  �E��E�    �M��E�    P�.{  j�E܋�P�E�P�$���M��|  �D��M�Q���   � �Ѓ�^��]� ��������U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �z  j �E܋�P�E�P�v#�����M����)|  ��t3���D��M�Q���   �@8�Ѓ����D��E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    �z  j�E܋�P�E�P��"���M��{  �D��M�Q���   � �Ѓ�^��]� ���U���$SV�E��E�    ���E�    P�M��E��  �E�    �E�    �y  j �E܋�P�E�P�f"�����M����{  ��t3���D��M�Q���   �@8�Ѓ����D��E�P���   �	�у���^[��]����������U���$�EV�E��E��E�   P�M��E��  �E�    �E�    �	y  h�   �E܋�P�E�P��!���M��}z  �D��M�Q���   � �Ѓ�^��]� �������t��t��t3�ø   ���̡D�Q�@L�@L�Ѓ���������������̡D�Q�@L�@P�Ѓ����������������U��D��u�u�@L�uQ���  �Ѓ�]� ������������U��D��uQ�@L��  �Ѓ�]� ��U��D��uQ�@L���   �Ѓ�]� �̡D�Q�@L�@X�Ѓ����������������U��D��u�u�@L�uQ�@\�Ѓ�]� ���������������U��D���0�@LSV��@�Ћ؅�u^[��]� W�M�����u�E��E�    �E؍M�D��E�    �E�    �E�    �E�    �]Ћ@h]  �@0�СD���j j S���   �@�Ѕ���   �D�S�@L�@�Ћ�������   �d$ �D����   �΋R(�ҋ��uԍE�Ph�   �  ����tq�M��tj�D�j ���   ���   �ЋЅ�tO�D�V���   �ʋ@<�СD��M�Q���   ���   �Ѓ���t�D�V�@@�@�Ѓ������d����*�D�S�@@�@�СD��M�Q���   ���   �Ѓ�3ۍM��p  �M����_^��[��]� ������������̡D�Q�@L�@`�Ѓ���������������̡D�Q�@L�@d�Ѓ����������������U��D��uQ�@L�@h�Ѓ�]� ����̡D�Q�@L��D  �Ѓ������������̡D�Q�@L�@l�Ѓ����������������U��D��uQ�@L���   �Ѓ�]� �̡D��@L�@�����U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@L���   ��Y�������������̡D�Q�@L���   �Ѓ�������������U���u�D��u�u�@L�u�u���   Q�Ѓ�]� ������U��D��u�u�@L�uQ���   �Ѓ�]� ������������U���u�D��u�u�@L�uQ��   �Ѓ�]� ���������U��D��u�u�@L�uQ��   �Ѓ�]� ������������U��D��@L��H  ]�������������̡D��@L��L  ��U��D��@L��P  ]��������������U��D��@L��T  ]��������������U��D��@L��p  ]��������������U��D��@L��t  ]��������������U��D��@L���  ]��������������U��D��@L���  ]��������������U��D��@L���  ]�������������̡D��@L���  ��U��U$V�u�EhP�h0�h �h�R�u �q�u�Q�u�D����@L�$�u���   VQ�Ѓ�4^]�  �������̡D��@���   ��D��@���   ��U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D�V�u�@�6���   �Ѓ��    ^]������������U��D�V�@L�@�Ћ���u^]áD�j �u�u�@�uV��h  �Ѓ���u�D�V�@@�@�Ѓ�3���^]������������U��D�j �u�H�E�� P�u��h  �u�Ѓ�]�������U��D��@���   ]��������������U��D��@L���   ]��������������U���u �D��u�u�@�u�u���   �u�u�Ѓ�]����U��� �D�W��E��E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4�D�jP�QL�΋��   �ЋE��E�E�Ph=���u��>
  ������   �D��M�Q���   ���   �Ѓ��E�    �M��y  ��^��]���U��� �D�W��E��E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4�D�jP�QL�΋��   �ЋE��E�E�Ph<���u��	  ������   �D��M�Q���   ���   �Ѓ��E�    �M���   ��^��]���U��D��@L���   ]��������������U��D��@L���   ]�������������̡D��@L��  ��D��@L��@  ��U��M�]� �����U��M�u��P]�U��M�u�u��P]��������������U���u�M�u�u��u�P]�������̡D����   �AP���   ��Y��������U��D��uQ�@8�@D�Ѓ�]� ����̡D��@8�@<�����U��D�V�u�@8�6�@@�Ѓ��    ^]���������������U���u�D��u�u�@8�u�u�@�uQ�Ѓ�]� ������U���u�D��u�u�@8�u�u�@Q�Ѓ�]� ��������̡D��@8� ������U��D�V�u�@8�6�@�Ѓ��    ^]���������������U��D��u�u�@8�uQ�@�Ѓ�]� ���������������U��D��u�u�@8Q�@�Ѓ�]� �̡D�Q�@8�@�Ѓ����������������U��D��uQ�@8�@ �Ѓ�]� �����U���u�D��u�u�@8�u�u�@$Q�Ѓ�]� ���������U��D��u�u�@8Q�@(�Ѓ�]� ��U��D��u�u�@8�uQ�@,�Ѓ�]� ���������������U��D��u�u�@8�uQ�@�Ѓ�]� ���������������U��D��u�u�@8Q�@0�Ѓ�]� ��U��D��u�u�@8�uQ�@4�Ѓ�]� ���������������U��D��uQ�@8�@8�Ѓ�]� �����U��M�D��P�APP�A@P�A0P�A P�AP���   Q�u�Ѓ�]�������������̡D��@���   ��D��@���  ��U��D��@�@,]�����������������U��D��@���  ]��������������U��D�V�uV�H�I�ыD�V�I�I8�у���^]����̡D��@�@<�����U��D��@�@@]����������������̡D��@�@D����̡D��@�@H�����U��D��@�@L]�����������������U��D��@�@P]�����������������U��D��@��<  ]��������������U��D��@��,  ]��������������U���u�D��u�u�@�u�u���   h�6  �Ѓ�]�����U��D��@�@]�����������������U��D��M��� �@Q�@�СD��M�j j�hl��@Q�@�СD��M�Q�@�@�СD��M�Q�M�Q�@�@�СD��M��� �@�@<�ЋD�j�j��u�Q�M�P�BL�СD��M�Q�@�@�СD��M�Q�@�@�СD��M�Q�@�@�Ѓ���]����U��D��@���  ]��������������U��D��@��8  ]��������������U��D��M����@VWQ��  �ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]����U��D��M����@VWQ��  �ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]����U��D��@��x  ]��������������U��D��@��|  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@�@T]�����������������U��D��@�@X]�����������������U��D��@�@\]����������������̡D��@�@`�����U��D��@���  ]�������������̡D��@�@d����̡D��@�@h�����U��D��@�@l]�����������������U��D��@�@p]�����������������U��D��@�@t]�����������������U��D��@��D  ]��������������U��D��@��  ]��������������U��D��@�@x]�����������������U��D��@��@  ]��������������U��V�u���"����D�V�u�I�I|�у���^]���������U��D��@���   ]��������������U��D��@��d  ]��������������U��D��@��h  ]��������������U��D��@���  ]�������������̡D��@���   ��U��V�u���R���D�V�I���   �у���^]��������̡D��@��`  ��U��D��@��  ]��������������U��D��M���@�uQ���   �ЋM���o ��~@��f�A��]������U��D��@���  ]��������������U���u�D��E���@�D$�E�$�u���   �Ѓ�]�����������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@��   ]��������������U��D��@��  ]��������������U��D��@��l  ]�������������̡D��@���  ��U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��M����@VW�u���  Q�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]�U��D��M����@VW�u���  Q�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]�U��D��@���  ]��������������U��D��@���  ]��������������U����D��U�R�U�R�@�U�RQ���   �Ѓ����#E���]����������������U����D��U�R�U�R�@�U�RQ���   �Ѓ����#E���]����������������U����D��U�R�U�R�@�U�RQ���   �Ѓ����#E���]����������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@���   ]��������������U��D��@��  ]��������������U��D��@��\  ]��������������U��D����u�H�E��uP��t  �у����v����M�������E��]��������U��D��@��H  ]��������������U��D��@��T  ]�������������̡D��@��p  ��U��D��@��8  ]��������������U���  ��3ŉE��EP�u������h   P��J ����x	=�  |#��D�h(�hH  �@��0  �Ѓ��E� �D�������Qhp��@��4  �ЋM���3��k�  ��]������������������������U���u(�E�u$�u �P�u�D��u�u�@0�u�u���   RQ�Ѓ�(]�$ ������U���u(�E�u$�u �P�u�D��u�u�@0�u�u���   RQ�Ѓ�(]�$ ������U���u(�D��u$�u �@0�u�u���   �u�u�u�uQ�Ѓ�(]�$ ���������̡D�Q�@0���   �Ѓ�������������U��D��u�u�@0Q���   �Ѓ�]� ���������������U���u�D��u�u�@0�uQ���   �Ѓ�]� ��������̡D�Q�@0���   �Ѓ�������������U���u�D��u�u�@0�uQ���   �Ѓ�]� ��������̡D��@0���   ��U��D�V�u�@0�6���   �Ѓ��    ^]������������U��D��M����@V�u�u��X  �uQ�Ћuj PV�    �F    �D����   �I�ыD��E�P���   �	�у� ��^��]����������U���4VhLGOg�M�����D�j P�E��IhicMCP��X  �ЋD����E�    �E�    j ���   �M�RQ�@�СD��M�Q���   � �Ѓ� �M��i���D��M�Q���   �@T�Ѓ���u
�M����� �D��M�Q���   �@T�ЋM��P����D��E�P���   �	�ыE��^��]������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��M����@VWj �u��t  �u�u�uQ�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у�(��_^��]������U��D��M����@V�u�u���  �u�uQ�Ћuj PV�    �F    �D����   �I�ыD��E�P���   �	�у�$��^��]�������U��D���4�@��p  �Ѕ���   h���M��U ���D��M��uh���@�@4�СD��M��uh���@�@4�СD��M�j Q�M��@hicMCQ��X  �ЋD����E�    �E�    j ���   �M�RQ�@�СD��M�Q���   � �СD��M�Q���   � �Ѓ�$�M��������]����������U��D���4�@V��p  �Ѕ�u�D��uV�H�I�у���^��]�Wh!���M��\����D��M��uh!���@�@4�СD��M�j Q�M��@hicMCQ��X  �ЋD����E�    �E�    j ���   �M�RQ�@�СD��M�Q���   � �СD��M�Q���   �@H�ЋD����}W�I�I�ыD�WV�A�@�ЋD��E�P���   �	�у�4�M��������_^��]������������U��D���4�@V��p  �Ѕ�u�D��uV�H�I�у���^��]�Wh����M��<����D��M��uh����@�@4�СD��M�j Q�M��@hicMCQ��X  �ЋD����E�    �E�    j ���   �M�RQ�@�СD��M�Q���   � �СD��M�Q���   �@H�ЋD����}W�I�I�ыD�WV�A�@�ЋD��E�P���   �	�у�4�M�������_^��]������������U��D���4�@��p  �Ѕ�u��]�Vh#���M��4����D��M��uh#���@�@4�СD��M�j Q�M��@hicMCQ��X  �ЋD����E�    �E�    j ���   �M�RQ�@�СD��M�Q���   � �СD��M�Q���   �@8�ЋD����E�P���   �	�у�(�M��������^��]�������U��D���4�@��p  �Ѕ�u��]�Vhs���M��T����D��M��uhs���@�@4�СD��M�j Q�M��@hicMCQ��X  �ЋD����E�    �E�    j ���   �M�RQ�@�СD��M�Q���   � �СD��M�Q���   �@8�ЋD����E�P���   �	�у�(�M��������^��]�������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@��@  ]��������������U��V�u���t�D�Q�@��D  �Ѓ��    ^]�������U��D��@��H  ]��������������U��D��@��L  ]��������������U��D��@��P  ]��������������U��D��@��T  ]��������������U��D��@��X  ]��������������U��D��@��\  ]�������������̡D��@��d  ��U��D��@��h  ]��������������U��D��@��l  ]��������������U��D��@���  ]�������������̡D��@���  ��U��D��@���  ]�������������̡D��@��P  ��D��@���  ��U��D��M���@�uQ���  �ЋM��P�����M������E��]���������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@��l  ]��������������U��D��@���  ]��������������U��D��@���  ]��������������U��D��@��$  ]��������������U��D��@��(  ]��������������U��D��@��,  ]�������������̡D��@��0  ��D��@��<  ��U��D��@��  ]��������������U��D��@��`  ]��������������U��D��@��\  ]��������������U��D��u�u�@TQ�@�Ѓ�]� ��U��D��uQ�@T�@�Ѓ�]� �����U��D��uQ�@T�@�Ѓ�]� �����U��D����u�@TQ�M�Q�@<�ЋM���o ��~@��f�A��]� �����U��D��@T� ]��U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�hG  �@T� �Ѓ�������������U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��D����E�@H�$Q�@�Ѓ�]� ����������̡D�j Q�@H���   �Ѓ�����������U��D��uj �@HQ���   �Ѓ�]� �D�jQ�@H���   �Ѓ�����������U��D��uj�@HQ���   �Ѓ�]� �D�jQ�@H���   �Ѓ����������U��D��uj�@HQ���   �Ѓ�]� �D�Q�@H���  �Ѓ�������������U��D��uQ�@H���  �Ѓ�]� ��U��D��uQ�@H���  �Ѓ�]� ��U��D��uQ�@H���  �Ѓ�]� ��U��D��u�u�@HQ��  �Ѓ�]� ���������������U��D��u�u�@HQ��  �Ѓ�]� ��������������̡D�Q�@H���   �Ѓ�������������U��VW�u���1�  ������t�D��uV�AHW���   �Ѓ���_^]� �������U��VW�u���u辊  ������t�D��uV�AHW���   �Ѓ���_^]� ����U��D��u�u�@HQ���   �Ѓ�]� ���������������U��D��u�u�@HQ���   �Ѓ�]� ���������������U��D��uQ�@H���   �Ѓ�]� �̡D�Q�@H���  �Ѓ�������������U���u�D��u�u�@H�u�u���  Q�Ѓ�]� ������U��D����@HWj �����   h�  W�Ѓ��} u�   _��]� Vh�  诈  ��������   �D�j VW�IH���   �у��M��R����D��M��uh�  �@�@0�СD��M��E���@�$h�  �@,�СD��M�j QV�@@�@(�Ѓ��M��Y���^�   _��]� ^3�_��]� �̡D�Q�@H���   ��Y��������������U��D��uQ�@H���  �Ѓ�]� ��U��D��uQ�@H���  �Ѓ�]� �̡D�Q�@H��4  �Ѓ�������������U��D��@H� ]��U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��S�]V�uW�; ���
  �D��uW�@H���   �Ѓ�����   �D�jW�@H���   �Ѓ�����   ��D�W�@H���   �Ѓ��} u!�u�D�S�u�@HV�u���  W�Ѓ��>��t:�u�D�S�u�@HV�u���  W�СD����΋��   �@(�Ћ���uɋu�; uS�D�W�@H���   �Ѓ���t;�    �D�W�@H���   �СD��uW�@H���   �Ѓ�_^[]� �   �   �D�W�@H���   �СD����} �@Hu!�u���  j �uV�uW�Ѓ���_^[]� � h  �Ћ؃���u_^[]� �D��΋��   �@x�ЋD�P���   �ˋB|�Ѕ�tP�u�D�j �u�@HV�u���  W�Ћȃ���t�D�S���   �@H�СD��΋��   �@(�Ћ���u�_^��[]� ����U���u�D��u�u�@H�u�u���  Q�Ѓ�]� �����̡D�Q�@H���   ��Y�������������̡D�Q�@H���   �Ѓ�������������U��D��u�u�@HQ���   �Ѓ�]� ��������������̡D�Q�@H���   ��Y�������������̡D�Q�@H��t  ��Y�������������̡D�Q�@H��P  �Ѓ������������̡D�Q�@H��T  �Ѓ������������̡D�Q�@H��X  �Ѓ�������������U��D����@HQ�M�Q��\  �ЋM���o ��~@��f�A��]� ����̡D�Q�@H��`  �Ѓ�������������U��D��uQ�@H��d  �Ѓ�]� ��U��D����E�@H�$Q��h  �Ѓ�]� ��������U��D����E�@H�$Q��t  �Ѓ�]� ��������U��D����E�@H�$Q��l  �Ѓ�]� ��������U��D��uQ�@H��p  �Ѓ�]� ��U���u�D��u�u�@H�uQ���  �Ѓ�]� ���������U���u�D��u�u�@H�u�u���  �uQ�Ѓ�]� ��̡D�h�  �@H� �Ѓ�������������U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@H���   �Ѓ������������̡D�Q�@H���   �Ѓ�������������U��D��uQ�@H���   �Ѓ�]� ��U��D��uQ�@H���   �Ѓ�]� ��U��D��u�u�@HQ���  �Ѓ�]� ���������������U��D��u�u�@HQ��   �Ѓ�]� ���������������U��D��u�E���@H�$���  Q�Ѓ�]� �����U��D�Vh  �@H� �Ћ�������   �uh�  豁  �Ѓ���t^�D�j RV�AH���   ���uh(  膁  �Ѓ���t3�D�j RV�AH���   �СD����΋��   j j�@�Ћ�^]áD�V�@@�@�Ѓ�3�^]�����U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@H��  �Ѓ������������̡D�Q�@H��  �Ѓ������������̡D�Q�@H���  �Ѓ������������̡D�Q�@H���  �Ѓ������������̡D�Q�@H���  �Ѓ�������������U��D��u�u�@HQ��  �Ѓ�]� ���������������U��D��u�u�@H�uQ��   �Ѓ�]� ������������U���u�D��u�u�@H�uQ��|  �Ѓ�]� ���������U��EV���u�D��@H���  �'��u�D��@H���  ���u(�D��@H���  V�Ѓ���tP�u���   ^]� 3�^]� ����������U���SW���  �؅���   �} ��   �D�Vj h�  �AHW��p  �ЋD���h�  W�u�IH���   �������E����   �u3��Ή}��  ����   �E���P�E�P�u�W��  ��t\�u�;u�T������u�U����ɋD�;D�t-�D��Hl����P�E�p�A�Ѓ��D����tP����  F;u�~��}��MG�}��  �u;��v���^_��[��]� _3�[��]� U����D�Vj ��@Hh�  V�u�p  �Ѓ��E���u^��]� �EW��u�D��@H���  �+��u�D��@H���  ����T  �D��@H���  V�Ћ������6  S���_  �D�3�h�  V�]��@H���   �Ѓ�����   �E��s���E�D��MS�@l�q�@�Ћ؃�����   �D��s�u�I\�I,�у���t�F���P�  �D��s�u�@\�@,�Ѓ���t�F���P�a  �M�;At"�D��s�u�@\�@,�Ѓ���tV���5  �D��s�u�@\�@,�Ѓ���t�F��P�  �D����]��ECh�  �@H�u�]����   �Ѓ�;�����[_�   ^��]� _3�^��]� ������̡D�Q�@H���  �Ѓ�������������U��D��u�u�@HQ���  �Ѓ�]� ���������������U��D��u�u�@H�uQ���  �Ѓ�]� �����������̡D�Q�@H���  �Ѓ������������̡D�Q�@H���  �Ѓ�������������U��D��uQ�@H��  �Ѓ�]� ��U��D��uQ�@H��  �Ѓ�]� �̡D�Q�@H��  �Ѓ�������������U��D��uQ�@H��  �Ѓ�]� �̡D�Q�@H��T  �Ѓ�������������U��D��u�u�@HQ��  �Ѓ�]� ���������������U��D��uQ�@H��8  �Ѓ�]� ��U��D��uQ�@H��<  �Ѓ�]� ��U��D��u�u�@H�uQ��@  �Ѓ�]� ������������U��D��uQ�@H���  �Ѓ�]� ��U��D��uQ�@H��H  �Ѓ�]� �̡D�Q�@H��L  ��Y��������������U��D�Vh�  �@H� �Ћ�����u^]áD��u�u�@HV��  �Ѓ���u�D�V�@@�@�Ѓ�3���^]����������U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��D��u�u�@H�uQ��   �Ѓ�]� ������������U��D����E�@H�$Q��$  �Ѓ�]� �������̡D�Q�@H��(  �Ѓ�������������U��D��u�u�@HQ��,  �Ѓ�]� ��������������̡D��@H��  ��U��D��@H��  ]�������������̡D�V��W�@@V�@,�ЋD����ȋBj h�  ���   �ЋD���h�  V�IH���   �у���
��t_3�^Ë�_^�̡D�Q�@@�@,�ЋD����ЋA��j h�  ���   �����U��D����E�u�@H�u����  �$Q�M�Q�ЋM���o ��~@��f�A��]� ��U��D����E�u�@H�u����  �$Q�M�Q�ЋM���o ��~@��f�A��]� �̡D�Q�@H���  �Ѓ�������������U��D��u�u�@HQ��8  �Ѓ�]� ���������������U���u�D��E���@H�$�u��0  Q�Ѓ�]� ��U��D��@H�@]�����������������U��D�V�u�@@�6�@�Ѓ��    ^]���������������U���u �D��u�E���@H�$�u���   �u�u�Ѓ�]�������������U���u�D��E���@H�$�u�u���   �u�Ѓ�]�����������������    ���������̡D�j�1�@H��|  �Ѓ����������U��D�V�u��@H��x  ��3ɉ��������^]� ���̡D�j �1�@H��|  �Ѓ����������U��fnE�M����YE�Xp��,�;�}��]�;EOE]����������������U���D�D�SVW�@H�}h�  W���   �ЋD�3�V��h�  �IHW�]Ћ��   �у��E��u�u��u���4	  �D��ϋ��   �@��=�  �D��n  �@HVh:  W���   �ЋD�h�  W�E�IH���   �ыD�Vh�  W�IH�E��uԋ��   �ыD���W�]�IH��  �ыD�W�E̋IH���  �у�(�E�3�9u���   �C3ۉE���$    �M̅�tNj�W��  ���t>�Mȍ@�|� ���M�~�� ��%�������;�u+��  �M�;�O��B�  ���E��M�� ;Au������E�G���E�;}�|��]ԋ]�E�}��tyj W���y  ���  �M��@y  ��t[�M��$s  �M�;�uL�D��Ih����h�  �@Q�M����  �Ѓ��EĉE����  �M���x  �u�P�u��$�  ���E�h��h�  �@�D���Q�M��@���  �Ѓ��E����}  �u��u�P��  �Mԃ���~,�D�h����h�  �@Q���   �Ѓ��E���;  �D�j�VW�@H��  �Ѓ����  �u��t jW���zx  ���  ���Kx  ���E��3��uܡD�j h�  W�@H���   �ЉE�3�3��U����E�9E���  �{�}����    �M̅��  j�P���  ����  �Mȍ@�|� �4��u�~�� ��%�������9E��2  ���@�  3ۉE�3��E�    9^~{��������Шte�E��������������u����E�T��E�N�L��J�E�L��E�N�L��J�E�L��E�N�uĉL��J�E�L���C;^|�����  �Ǚ+�����~�M�QPQ�M���
  �U�3��]��M܍R�ÉE��+ÉEċƍI ;E���  �E����t.�E�[�oȋM�E���E�[�~D��E�M�f�D�E��[�oȋM���[�~D��M�f�A;�}j�E�9�u_�L�������������w>�$�x��M���U����-�M���U��T���M���U��T���M���U��T���U���;�|��M�E؃�B�M�M�@�U��E�;�����;E���  �}��_  �U��3�;G�M��Å���   �R�ƋG��@�o���~D�f�B�G��@�E��o��B�~D�f�B(��U��@�E�ȍR�o�D�0�~Af�D�@��t%�G�@�E��oȍȍR�D�H�~Af�D�X�G��u��@�E��oȍȍR���~Af�D��G��W�B�@�E��oȍȍR���~Af�D���W�B�@�E��oȍȍR���~Af�D��B�U���t-�G�@�E��oȍȍR���~Af�D��WB�U����G��}ЋU��Eԃ��u�@�Eԉ}�;E��i����E�P�0����E�P�'������  �E�P�����E�P�����E�P������3�_^[��]Ë��   �ϋ@��=  ��  �D�j h(  W�@H���   �ЋD���h(  W�IH���   �у��E�3Ʌ�~�I �˅�t�|� �4Vu���A;�|�E�h��hY  �@�D���Q�M��@���  �Ѓ��E�����   �u��u�P薳  �E�h��h^  ��    �D�Q�M��@���  �Ѓ��E��tD�u�SP�Z�  �D��ƙ+����IHPVW��   �E��у���u�E�P�ܯ���E�P�ӯ����_^3�[��]áD�j h�  W�@H���   �ЋD�j h(  W�IH�E����   �ы�3��E�3ۃ��M�3҉u��]؅���   �}䐋߅���   3��EЃ�~d�M��X�R�4v�����E��I0�EЍvC���oD��A��~D�f�A��E��o�A��~D�E�f�A��}�;ǋE�|��u��]؃|� tL�}�ƍ@�E��oȍȍRB���~A�vf�D��E��oȍȍRB���~Af�D��}�4ߋEԉu�C�]�;������MċU�3���~�I �D�    ��   @;�|�E�P�c������E�P�W�����_^�   [��]Þ���������������U���u�D��E���@H�$�u�u���  �Ѓ�]���U��D��@H���  ]��������������U��D��@H���  ]��������������U���u0�E(�D����@H�$�u$�u ���  �u�u�u�u�u�u�Ѓ�,]�U��D��@H���  ]��������������U��D��@H���  ]��������������U���u0�E�u,�D��u(�u$�@H�u ����P  �D$�E�$�u�u�Ѓ�,]������������������A    ��q����D��@l�@��Y���������U��D�V��@l�v�@�ЋM����u�A^]� �D��u�u�@lQ�u� ��3ɉF��������^]� �������������̋I��u3�áD�Q�@l�@�Ѓ������U����D��U�R�U�R�u�@l�u�q�@�ЋM����U;�u	�E���]� ���9U�D���]� �������U��D��@H���   ]��������������U��D��@H���  ]��������������U����D����MW��@�$�u���   ���E�]��M�f/�w�Ef/�w(��D����M�@�$�u�@,�Ћ�]����������U���H�D��M�W�Q�ufE�M��E��@Q�M���   ���M�o �~`�E��Ef/�v(��	f/�v(��U�f/�v(��	f/�v(��]�f/�wf/�v(��(áD��M��E��U��e��@Q�u�M�@H�Ћ�]��������U��D��@H��0  ]�������������̋������������������������������̡D��@H���  ��U��D��@H���  ]��������������U���u0�D��u,�u(�@H�u$�u ���  �u�u�u�u�u�uQ�Ѓ�0]�, ����U���u0�D��u,�u(�@H�u$�u ���  �u�u�u�u�u�uQ�Ѓ�0]�, ���̡D�Q�@H��,  �Ѓ�������������U��D��uQ�@H��X  �Ѓ�]� �̡D�Q�@H��\  �Ѓ�������������U��D�Q�u�@H�u���   �Ѓ�]� ���������������U��QSV��3ҋM���u�W�}�σ�t
����B��u��PSWV�M�	  �} ~(��   VW�}��MW�o  SVW�M��  _^[��]� ;�tSWV�M�L  _^[��]� ���U��V���v����D��@l�@�Ѓ��Et	V�է������^]� �����������U���V�u����   �ƙ+U����AS�Z��M�W�	�<�E��ˉ}�]���d$ �]��}�E���$    ��~I�����M��]��E��*�G����N�S��G�C�u�}��W��~g�M��U����9u����    ���G���;�}��U;H}G���;�M��w������s��H�K�?�p�u��U;�~��M��N���_[^��]� �����U��UV�u��+����� ~^�E�U]�����S�ZW�]��I ��;�t7�]��$    �;H�}�p�ыH���H��H�P��p����;�u܋]�U�u���];�u�_[^]� ��U��Q�U��W�}+ǃ���M�=   ��   S�]V�E����   H�J��E��+����+���4Ǎǋ;�}
;�|��;��
;�}���;�Lًu�}������9|���    ��;|�;�s$���V��G�F��W;�u����;�uƋ����u�]�u�M�VS�>����}��+��U�����   �J���^[_��]� �M�RWS����^[_��]� ��������U��QS�]V�u;�t8W��F���;}$���N�M���@��
�R��H�J;8|�E��:�B��;�u�_^[��]� �D�Q�@\�@�Ѓ���������������̡D�Q�@\�@�Ѓ����������������U��D��uQ�@\�@�Ѓ�]� �����U��D��u�u�@\Q�@�Ѓ�]� ��U��D��uQ�@\�@�Ѓ�]� ����̡D�Q�@\�@�Ѓ����������������U��D��uQ�@\�@ �Ѓ�]� �����U��D��u�u�@\Q�@$�Ѓ�]� ��U���u�D��u�u�@\�uQ�@`�Ѓ�]� ������������U��D��uQ�@\�@0�Ѓ�]� �����U��D��uQ�@\�@@�Ѓ�]� �����U��D��uQ�@\�@D�Ѓ�]� �����U��D��uQ�@\�@H�Ѓ�]� ����̡D�Q�@\�@4�Ѓ����������������U��D��u�u�@\Q�@8�Ѓ�]� ��U��D��uQ�@\�@<�Ѓ�]� �����U���SVW�}��j �ω]�膻���D�S�@\�@�Ѓ��؋�S�k���3���~?��I �D��M�Q�MQ�@\h���V�u��@`�Ѓ����u�5����u����+���F;�|�_^[��]� �������������U���S�]�E�W����P舾���}� |z�D�W�@\�@�Ѓ��E���P�f����E���tWV3���~B�E��P�M����E���P�B����M;M��D�QW�@\�@�ЋM��A�M;M�~�F;u�|�^_�   [��]� _�   [��]� ����������̡D��@\� ������U��D�V�u�@\�6�@�Ѓ��    ^]��������������̸   � ��������3�� �����������3�� ����������̸   @� ��������3�� ����������̸   � ��������U��D��u�H�I�ыE��]� ��̸   � ��������U����   V�u��u3�^��]�h�   ��@���j P�Ū  �E�E��E�E��Eh�   ��@�����@���P�u��`����uǅD����j�E�#��E�-��E�s��E�2��E�X��E�n��E�(��E�7��϶���� ^��]��������U����   h�   ��@���j P�$�  �Eh�   �E���@���P�uǅ`���    �uj�{����� ��]�����U���   SV�u(3�W3��]����w  �D��M�@�@<�Ѕ��F  �����E�����   �EP�M�������D��M�Q�@�@�СD��M�Wj�h���@Q�@�Ѓ��E�M�P�š���u��E�Wj�P�E�P��\���P�_?������P��x���P�������P�E�P��������P�����E���t�E� �� t�M����������t��x�������С����t��\������轡����t�M̃��譡����t�D��M�Q����@�@�Ѓ���t�M�脡���}� t�u(�u$�u��u�u�u���������E�P�Y������V�u$j �u�u�u�p��������D��EP�I�I�у���_^[��]Ë�`��`��`��` ��`����U��M�EQj�u��E�A�Խ����]���������������̸   �����������U��V�u��t���u6j�u�ս������u3�^]Ë��B����ȅ�t��t��E3�;AOʋ�^]�������V���$��F    �D��@4���   �ЉF��^����������V���v�$��D��@4���   �Ѓ��F    �F    ^��� �������������U����u��U��u�E�    �u�E�    �u�uR�U�R�P�E�3Ɂ}�gnolE���]� �����������U���u�D��u�u�@4�u�u���   �u�q�Ѓ�]� ̡D��q�@4���   ��Y�����������̡D��q�@4���   ��Y������������U��D��u�q�@4���   �Ѓ�]� �D��q�@4���   �Ѓ�����������U���u�D��u�u�@4�q���   �Ѓ�]� ����������U���u�D��u�u�@4�q���   �Ѓ�]� ����������U��EQh`�u�P�D�R�q�@4���   �Ѓ�]� ���U��D��u�u�@4�q���   �Ѓ�]� �������������V���$��F    �D��@4���   �Ћ��0��V�D�R�A4���   �СD����@4���   �ЉF��^����������V���v�$��D��@4���   �Ѓ��F    �F    ^��U��D��u�u�@4�q���   �Ѓ�]� �������������U��D��u�u�@4�q���   �Ѓ�]� �������������U��D��u�u�@4�q���   �Ѓ�]� ������������̡D��q�@4���   �Ѓ�����������U���u�D��u�u�@4�q���   �Ѓ�]� ����������U��D��u�q�@4���   �Ѓ�]� U��D��u�q�@4���   �Ѓ�]� U��D��u�q�@4���   �Ѓ�]� U��D��u�q�@4���   �Ѓ�]� U��D��u�u�@4�q���   �Ѓ�]� �������������� �������������U��D��u�u�@4�q���   �Ѓ�]� �������������U��M��t�u$��u �u�u�u�u�u�P]�����������U��V���v�$��D��@4���   �Ѓ��F    �E�F    t	V�t�������^]� �����������    ���A    �A    �A    ���V��~ u=���t�D�Q�@<�@�Ѓ��    W�~��t������W�������F    _^���������U����E�VP���^�������P�   �M���ɚ����^��]���U��V��~ u1jh8�j;j��������t�u���S����3��F��u^]� �~ t3�9^��]� �D��u�@<� �Ћ��F   ���3�����^]� ��������V���F   �D��@<�@��3ɉ��^�����������������U��	�D���u	�@� ]� �@<�uQ�@�Ѓ�]� �����̃y t�   ËQ��u3�áD�R�1�@<�@�Ѓ��������V��~ u=���t�D�Q�@<�@�Ѓ��    W�~��t���{���W�u������F    _^���������U�����D���u�@� ]Ë@<�uQ�@�Ѓ�]�������U������$V��u�D��A�0��D��uQ�@<�@�ЋD������I�E�SP�I�ѡD��M�QV�@�@�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M��� �@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD�����[t(�H�uV�I�ыD��E�P�I�I�у���^��]Ë@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��uV�@�@�СD�V�H�E�P�I�ыD��E�P�I�I�у���^��]������������U������$SV��u�D��A�0��D��uQ�@<�@�ЋD������I�E�P�I�ѡD��M�QV�@�@�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M��� �@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD�����t)�H�uV�I�ыD��E�P�I�I�у���^[��]Ë@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD������?����@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��uV�@�@�СD�V�H�E�P�I�ыD��E�P�I�I�у���^[��]���U������$SV��u�D��A�0��D��uQ�@<�@�ЋD������I�E�P�I�ѡD��M�QV�@�@�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M��� �@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD�����t)�H�uV�I�ыD��E�P�I�I�у���^[��]Ë@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD������?����@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD�����������@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��uV�@�@�СD�V�H�E�P�I�ыD��E�P�I�I�у���^[��]�����������U������$SV��u�D��A�0��D��uQ�@<�@�ЋD������I�E�P�I�ѡD��M�QV�@�@�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M��� �@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD�����t)�H�uV�I�ыD��E�P�I�I�у���^[��]Ë@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD������?����@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD�����������@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��M�Q�@�@�СD��M�j j�h|��@Q�@�СD��M����@j Q�M܋@@Q�M��Ѕ��MܡD�Q�Ë@�@�СD����������@�M�j�u��@H�СD��M�j�j��u�@�u��@L�СD��uV�@�@�СD�V�H�E�P�I�ыD��E�P�I�I�у���^[��]���U��E�����EȉM]��  ������U��D��@<�@]�����������������U��E����u��]�VP�M��Չ���E�E�    P�E��E    P�M���������   �u�E���tA��t<��uX�D��u���   �@H�ЋD��Ѓ��A��V�@x�Ѕ�u+�   ^��]áD��u���   �@T��VP�Y�������uՍEP�E�P�M�肉����u�3�^��]��������U���DS3ۍM܉]��D�VQ�@�@�СD��M�Sj�h���@Q�@�СD��M�Q�@<�@�ЋD����E�P�I�I�у���u^3�[��]�WV�M�3�詈���E�P�E�P�M��������  ��}���   �D��u����   �@T�Ћ�������   �D����A�M�Q�@�СD��M̃��@Qj�M����   Q���ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M܃��@�u�@x���E���t�E� ��t�D��M�Q����@�@�Ѓ���t�D��M�Q����@�@�Ѓ��}� u!�E�P�E�P�M��ڇ�����������_^[��]Ë}���_^[��]��������������U���@SV�u3ۉ]���u^�D��M�Q�@�@�СD��M�Vj�h���@Q�@�СD��M�Q�@<�@�ЋD����E�P�I�I�у���u^3�[��]�V�M������E�P�E�P�M��%�����t�W�}�E�����   �D��u����   �@T�Ћ�������   �D����A�M�Q�@�СD��MЃ��@Qj�M����   Q���ЋD����E�P�I�I�ыD��A�M�QV�@�СD��M�Q�@�@�СD��M����@W�@x���E��t�E ��t�D��M�Q����@�@�Ѓ���t�D��M�Q����@�@�Ѓ��} tA�E�_^[��]Ã�u2�M���t+�D�Q���   �@H�ЋD��Ѓ��A��W�@x�Ѕ�t��E�P�E�P�M��օ���������_^[��]�������̡D��@<�@����̃=�� uK�����t�D�Q�@<�@�Ѓ����    V�5����t��� ���V���������    ^������������3�� �����������3�� �����������3��  ����������̸   � ��������3�� �����������3�� ���������������������������3�� �����������3�� ������������ �������������3�� �����������U���   ������h   j P�T�  �u �������u�u�u�uP�)   h   ������P�u�uj
蠝����8��]����������U��V�u�u�uj �u�uV赸���E�����   ǆ�   �ǆ�   �ǆ�   iǆ�   �ǆ�   �ǆ�   �ǆ�   ǆ�   �ǆ�   Uǆ�   �ǆ�   �^]Ë�`L��`\��``��`d��`h��`l���������̸   � ��������3�� �����������3�� ������������ �������������U��EW� �@]� �����������3�� �����������3�� ������������ �������������� �������������3�� �����������U��D���   �M�@�@<�Ѕ�tj �u�u�&�������u��]�h   ������j P�X�  �u �������u�u�uP�    h   ������P�u�uj觛����4��]�U��V�u�u�uj �u�uV�Ŷ����ǆ�   �ǆ�   �ǆ�   �ǆ�   iǆ�   Uǆ�   �ǆ�   �ǆ�   �ǆ�   �ǆ�   �^]Ë�`D��`H��`X������������U��Vj j�u����������t�@��t	����^]� 3�^]� U��Vj j�u���^�������t�@��t	����^]� 3�^]� U��Vj j�u���.�������t�@��t����^]� �������U��Vj j�u�����������t�@��t	����^]� 3�^]� U��Vj j�u�����������t�@��t	����^]� 3�^]� U��Vj j�u����������t�@��t	����^]� 3�^]� U��Vj j �u���n�������t�@ ��t�u����^]� 3�^]� �������������U���(Vj j$�u���+�������t^�@$��tW�M�Q���Ћu�Vj �����    �B    �D�PR���   �I�ыD��E�P���   �	�у���^��]� �D��M��E�    �E�    �E������E�    �E�    ���   j Q�M��@Q�СD��M�Q���   � �Ћu�E؍Vj ��    �B    �D����   �E�PR�I�ыD��E�P���   �	�у� ��^��]� �������U��Vj j(�u����������t�@(��t�u����^]� ����U��Vj j,�u�����������t�@,��t	����^]� 3�^]� U��Vj j0�u����������t�@0��t	����^]� 3�^]� U��E�@_�@b��@]��@Z�@g��@l��@ d�@$q��@(��@,i�@0��@4U]�����3�� ��`T��`(��`,��`<��`P��U��EVW�9�0;�t_3�^]� �P��u ��u9pu9qu��u�9yu�_�B^]� S�Y��u"��u9yu��u3��u/9pu*[_�   ^]� ��t��t;�u�P��t�A��t�;�t�[_3�^]� U���u�e������@]� ������������Vh��j\hD ���L�������t�@\��tV�Ѓ���^�����U��Vh��j\hD ����������t2�@\��t+V��h��jxhD ���������t�@x��t	V�u�Ѓ���^]� ���������U���Vh��j\hD ����������tG�@\��t@V�ЋEh��jdhD �E��E�    �E�    ��������t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��j\hD ���9�������t2�@\��t+V��h��jdhD ��������t�@d��t	�uV�Ѓ���^]� ���������U��Vh��j\hD �����������tZ�@\��tSV��h��jdhD ��������t�@d��t	�uV�Ѓ�h��jhhD ��������t�@h��t	�uV�Ѓ���^]� �U��Vh��j\hD ���Y���������   �@\��t{V��h��jdhD �3�������t�@d��t	�uV�Ѓ�h��jhhD ��������t�@h��t	�uV�Ѓ�h��jhhD ���������t�@h��t	�uV�Ѓ���^]� �����Vh��j`hD ����������t�@`��tV�Ѓ�^�������U��Vh��jdhD ���y�������t�@d��t	�uV�Ѓ�^]� �������������U��Vh��jhhD ���9�������t�@h��t	�uV�Ѓ�^]� �������������Vh��jlhD �����������t�@l��tV�Ѓ�^�������U��Vh��jphD �����������t�@p��t�uV�Ѓ�^]� ���^]� ���U��Vh��jxhD ����������t�@x��t	V�u�Ѓ���^]� �����������U��Vh��j|hD ���I�������t�@|��tV�u�Ѓ�^]� 3�^]� ������U��Vh��j|hD ���	�������t�@|��tV�u�Ѓ����@^]� �   ^]� ��������������U���Vh��jthD ����������tP�@t��tI�u�M�VQ�Ћu����P�`���h��j`hD ��������th�H`��ta�E�P�у���^��]� h��j\hD �N����u����t4�@\��t-V��h��jdhD �)�������t�@d��th��V�Ѓ���^��]� �������U��Vh��h�   hD �����������t���   ��t�uV�Ѓ�^]� 3�^]� U��Vh��h�   hD ����������t���   ��t�uV�Ѓ�^]� 3�^]� VW��3����$    �h��jphD �_�������t�@p��t	VW�Ѓ������8 tF��_��^�������U��SV��3�W��    h��jphD ��������t�@p��t	VS�Ѓ������8 tph��jphD ���������t�@p��tV�u�Ѓ�������h��jphD ��������t�@p��t	VS�Ѓ�����W���x�����tF�^����E_��t�0��~=h��jphD �_�������t�@p��t	VS�Ѓ������8 u^�   []� ^3�[]� �����������U���Vh��h�   hD ����������t<���   ��t2�u�M�VQ��h��j`hD ���������t�@`��t	�M�Q�Ѓ���^��]� �������U���Vh��h�   hD ��������tS���   ��tI�u�M��uQ�Ћu����P�:���h��j`hD �Y�������td�H`��t]�E�P�у���^��]�h��j\hD �*����u����t2�@\��t+V��h��jxhD ��������t�@x��t	V�u�Ѓ���^��]�������̋���������������h��jhD ��������t	�@��t��3��������������U��V�u�> t+h��jhD ��������t�@��tV�Ѓ��    ^]�������U��} W��t0h��jhD �C�������t�@��t�u�uW�Ѓ�_]� 3�_]� �������������U��Vh��jhD �����������t�@��t�uV�Ѓ�^]� 3�^]� ������U��Vh��jhD ����������t�@��t�uV�Ѓ�^]� 3�^]� ������Vh��j hD ���|�������t�@ ��tV�Ѓ�^�3�^���Vh��j$hD ���L�������t�@$��tV�Ѓ�^�3�^���U��Vh��j(hD ����������t�@(��t�u�u�uV�Ѓ�^]� 3�^]� U��Vh��j,hD �����������t�@,��t�u�uV�Ѓ�^]� 3�^]� ���U��Vh��j(hD ����������t�@0��t�u�u�uV�Ѓ�^]� 3�^]� Vh��j4hD ���\�������t�@4��tV�Ѓ�^�3�^���U��Vh��j8hD ���)�������t�@8��t�u�u�u�uV�Ѓ�^]� 3�^]� �������������U��Vh��j<hD �����������t�@<��t	�uV�Ѓ�^]� �������������U��Vh��h�   hD ����������u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ���V�������u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ����������u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD �����������t�u���   �u�uV�Ѓ�^]� �����Vh��jDhD ����������t�@D��tV�Ѓ�^�3�^���U��Vh��jHhD ���i�������t�u�@HV�Ѓ�^]� �U��Vh��jLhD ���9�������u^]� �u�@LV�Ѓ�^]� ������������U��Vh��jPhD �����������u^]� �u�@P�uV�Ѓ�^]� ���������U��Vh��h�   hD ����������u^]� �u���   �u�uV�Ѓ�^]� U��Vh��h�   hD ���v�������u^]� �u���   �u�u�u�uV�Ѓ�^]� ����������Vh��jThD ���,�������u^Ë@TV�Ѓ�^���������U��Vh��jXhD �����������t�u�@XV�Ѓ�^]� �U���Vh��h�   hD �����������tQ���   ��tG�u�M�Q���Ћu��P�l���h��j`hD ��������t|�H`��tu�E�P�у���^��]� h��j\hD �E�    �E�    �E�    �E����u����t3�@\��t,V��h��jdhD � �������t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��h�   hD �����������t���   ��t�u���u�u��^]� 3�^]� ������������U��Vh��h�   hD ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   hD ���F�������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   hD ����������t���   ��t�u����^]� 3�^]� ��Vh��h�   hD �����������t���   ��t��^��3�^����������������U��Vh��h�   hD ����������t���   ��t�u���u�u��^]� 3�^]� ������������U��Vh��h�   hD ���6�������t���   ��t�u����^]� ���������U��Vh��h�   hD �����������t���   ��t�u���u�u��^]� 3�^]� ������������Vh��h�   hD ����������t���   ��t��^��3�^����������������U��h��jhD �l�������t
�@��t]��3�]��������U���Vh��h�   hD �5�������u�D��uV�H�I�у���^��]Ë��   �M�W�uQ�ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]���U��h���uhD ������]�������Vh��h�   h D ����������t���   ��t��^��3�^����������������Vh��h�   h D ���I�������t���   ��t��^��3�^����������������Vh��h�   h D ���	�������t���   ��t��^��^��U��Vh��h�   h D �����������t���   ��t�u����^]� 3�^]� ��Vh��h�   h D ����������t���   ��t��^��^��U���Vh��h�   h D ���c�������t=���   ��t3�E�M���$Q���ЋM^�o ��~@��f�A��]� �EW�^ �@��]� ����������Vh��h�   h D �����������t���   ��t��^��3�^����������������U��Vh��h�   h D ����������t���   ��t�u����^]� ���^]� �U��Vh��h�   h D ���f�������t���   ��t�u����^]� 3�^]� ��U���8Vh��h�   h D ���#�������tG���   ��t=�u�M�Q���ЋM^�o ��o@�A�o@ �A �~@0��f�A0��]� �EW�( ����^�@0    � ���f�H�H�P �@(��]� ���������������U��Vh��h�   h D ���f�������t���   ��t
�u���u��^]� ������U���Vh��h�   h D ���#�������tZ���   ��tP�u�M�Q���Ћuj PV�    �F    �D����   �I�ыD��E�P���   �	�у���^��]� �E^�     �@    ��]� �����������U��Vh��h�   h D ����������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h D ���6�������t���   ��t�u����^]� 3�^]� ��Vh��h�   h D �����������t���   ��t��^��3�^����������������Vh��h�   h D ����������t���   ��t��^��3�^����������������Vh��h�   h D ���y�������t���   ��t��^��3�^����������������Vh��h�   h D ���9�������t���   ��t��^��3�^����������������Vh��h�   h D �����������t���   ��t��^��^��U��MVh!D �u�܏������t+h��h�   h D ��������t���   ��t��^]��^]���������h��h�   h D �|�������t���   ��t��3��������U��h��h�   h D �I�������t���   ��tV�u�6�Ѓ��    ^]ËE�     ]����������Vh��h�   h D �����������t���   ��t��^��3�^����������������U��Vh��h�   h D ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h D ���v�������t���   ��t�u����^]� ���^]� �U��Vh��h�   h D ���6�������t���   ��t
�u���u��^]� ������U��h���uh D �������]�������U��U�f.���D��   �Af.B���D��   �Af.B���Dzy�A;Buq�A f.B ���Dza�A(f.B(���DzQ�A0f.B0���DzA�A8f.B8���Dz1�A@f.B@���Dz!�AHf.BH���Dz�A;Bu	�   ]� 3�]� �����U���u�5������@]� ������������h,�h  h�e ���������t��  ��t��3��������U��h,�h  h�e ���������t��  ��t]��]����Vh,�h�   h�e ����������t���   ��t��^�����^���������������U��Vh,�h�   h�e ���V�������t���   ��t�u����^]� 3�^]� ��U���Vh,�h�   h�e ����������t=���   ��t3�E�M���$Q���ЋM^�o ��~@��f�A��]� �EW�^ �@��]� ����������Vh,�h�   h�e ����������t���   ��t��^��^��U��Vh,�h�   h�e ���f�������t���   ��t�u����^]� 3�^]� ��U��Vh,�h$  h�e ���&�������t��$  ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e �����������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ����������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ���f�������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ���&�������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e �����������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ����������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ���f�������t���   ��t�u����^]� 3�^]� ��U��Vh,�h  h�e ���&�������t��  ��t�u���u��^]� 3�^]� ���������������Vh,�h  h�e �����������t��  ��t��^��^��Vh,�h�   h�e ����������t���   ��t��^��^��Vh,�h�   h�e ���y�������t���   ��t��^��^��Vh,�h�   h�e ���I�������t���   ��t��^��^��Vh,�h�   h�e ����������t���   ��t��^��^��U��Vh,�h  h�e �����������t��  ��t�u���u��^]� 3�^]� ���������������U��Vh,�h   h�e ����������t��   ��t�u���u��^]� 3�^]� ���������������U��Vh,�h<  h�e ���F�������t��<  ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ����������t���   ��t�u����^]� ���������Vh,�h�   h�e �����������t���   ��t��^��3�^����������������U��Vh,�h  h�e ����������t%��  ��t�u���u�u�u�u�u��^]� 3�^]� ���U��Vh,�h  h�e ���6�������tR��  ��tH�E0��0���D$(�E(�D$ �E �D$�E�D$�E�D$�E�$��^]�0 ��������U��Vh,�h(  h�e ��趿������tR��(  ��tH�E0��0���D$(�E(�D$ �E �D$�E�D$�E�D$�E�$��^]�0 ��������U��Vh,�h�   h�e ���6�������t.���   ��t$�u�E�΃��D$�E�$��^]� ���^]� ���������U��Vh,�h�   h�e ���־������t���   ��t�u����^]� 3�^]� ��U��Vh,�h0  h�e ��薾������t��0  ��t�u����^]� 3�^]� ��U��Vh,�h,  h�e ���V�������t��,  ��t
�u���u��^]� ������U��Vh,�hD  h�e ����������t��D  ��t�u����^]� 3�^]� ��U��VWh,�h�   h�e ���ս��������tG���    t>j<j h���e  ����� C���0C�ϋ��   �uh(�j<h����_^]� ���������������Vh,�h�   h�e ���Y�������t���   ��t��^��3�^����������������U��Vh,�h�   h�e ����������t���   ��t�u����^]� 3�^]� ��U��Vh,�h�   h�e ���ּ������t���   ��t�u����^]� ���������U��Vh,�h�   h�e ��薼������t���   ��t�u����^]� ���������Vh,�h�   h�e ���Y�������t���   ��t��^��3�^����������������Vh,�h�   h�e ����������t���   ��t��^��3�^����������������U��Vh,�h   h�e ���ֻ������t ��   ��t�u���u�u�u�u�u��^]� ����������U��Vh,�h@  h�e ��膻������t)��@  ��t�oE���΋��u� �~Ef�@��^]� �U��Vh,�h4  h�e ���6�������t��4  ��t�u���u�u��^]� ���U��Vh,�h8  h�e �����������t��8  ��t�u���u�u��^]� ���U��Vh,�hH  h�e ��趺������t��H  ��t�u���u��^]� 3�^]� ���������������U��M���E��D$�E�$�]� ����������U��M���E��D$�E�$�u�P]� ������U��h,��uh�e ������]�������U��h0�jhD ��������t
�@��t]��3�]��������U��h0�jhD 輹������t
�@��t]��]����������U��h0�j8hD 茹������t
�@8��t]��]����������U��QVh0�j8hD �Z���������th�~8 tb�D����   ���   �ЉE���t-�D��u���   �ȋ��   ���u�F8�u�u��u�Ѓ��D��M�Q���   ���   �Ѓ�^��]�����h0�jhD �ϸ������t	�@��t�����������������U��h0�jhD 蜸������t
�@��t]��3�]��������U��V�u��u3�^]áD����   ���   �ЉE��tF�D�V���   �ȋ��   �Ћuh0�jhD �+�������t�@��t�uV�Ѓ����3��D��MQ���   ���   �Ѓ���^]����������������U��h0�j4hD �̷������t
�@4��t]��3�]��������U��h0�j hD 蜷������t
�@ ��t]��3�]��������U��h0�j$hD �l�������t
�@$��t]��3�]��������h0�j(hD �?�������t	�@(��t��3��������������U��h0�j,hD ��������t
�@,��t]��3�]��������h0�j0hD �߶������t	�@0��t��3��������������U��h0��uhD 諶����]�������h4�jhD 菶������t	�@��t��3��������������U��h4�jhD �\�������t
�@��t]��3�]��������U����o���D����u�u�A�ʋ��   �ЋE��B����} tj�%n����]� j �n����]� U��U��3ɋ���tvV�u;�t�D�A���u�^��]� �D����tS�E�   �E��=o���D��ЋA�M�Q�u�ʋ��   �СD��M�Q���   � �ЋE�裀��j �m����^��]� ��U����n���D����u�A�ʋ@t�ЋD�j P�u���   �A�ЋE���]� ���������������U���V�n���D����u�A�ʋ@t�ЋD�P���   �@8�ЋU����3��:�tZ��9qt@�<����u�^��]� �M��E��D��E�   j Q���   �u�@�СD��M�Q���   � �ЋE���^��]� �������������U���V�u�E�    W����   �}��u��m�����D��E�    �E�    S�A�ϋ]S�@t�ЋD��Ћ��   �M�QR�@�Ѓ���uC�D���S�@�@t�ЋD�P���   �@�ЋD����u���   �I�у�;�u2����D��M�Q���   � �Ѓ���[td�D����u�u�@���   ��_^��]� ���/����}��tj P���.�����t(j W���`����Ѕ�t�D��uj�A�ʋ��   ��_^��]� ����������V���hN�������^���������������U��V�uj �u�uj �uV��   ����u3�^]�j#V��N��������t�D�V�@@�@,�ЋD����ЋA���uh�  �@4�СD�V�@@�@,�ЋD����ЋA���uh�  �@4�Ћ�^]���������������U��h4��uhD �K�����]�������U��V�uW�u�}j W�u�uV�Á�������   _^]�������U��D���   �@V�u�΋@<�Ѕ�tj V�u�u�������u^��]�h   ������j P�Y  �u������j j V�u�uP�L���h   �������u�P�u�uj#��e����8^��]���������Vh8�jh�t����l�������t�@��t��^��3�^������Vh8�jh�t����<�������t�@��t��^��3�^������U���Vh8�jh�t�����������tV�@��tOW�u�M�Q���ЋD����}W�I�I�ыD�WV�I�I�ыD��E�P�I�I�у���_^��]� �D��uV�H�I�у���^��]� ������������Vh8�jh�t����l�������t�@��t��^��3�^������U��Vh8�jh�t����9�������t�@��t�u���u��^]� 3�^]� �����U��Vh8�j h�t������������t�@ ��t�u���u��^]� 3�^]� �����Vh8�jh�t���輯������u^Ë@V�Ѓ�^���������U��h8��uh�t�苯����]�������U��Vh@�h�   h�f ���f�������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh@�h�   h�f ����������t���   ��t�u���u��^]� ���^]� ��������������U��Vh@�h�   h�f ���Ʈ������t���   ��t�u����^]� 3�^]� ��U��Vh@�h�   h�f ��膮������t���   ��t
�u���u��^]� ������U��Vh@�h�   h�f ���F�������t���   ��t�u����^]� 3�^]� ��U��Vh@�h�   h�f ����������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh@�h�   h�f ��趭������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh@�h�   h�f ���f�������t���   ��t�u����^]� 3�^]� ��Vh@�h�   h�f ���)�������t���   ��t��^��3�^����������������U��Vh@�h�   h�f ����������t���   ��t�u����^]� 3�^]� ��U��Vh@�h�   h�f ��覬������t���   ��t�u���u��^]� 3�^]� ���������������Vh@�h�   h�f ���Y�������t���   ��t��^��3�^����������������U��Vh@�h�   h�f ����������t���   ��t�u����^]� 3�^]� ��U��V�u�> t2h@�h�   h�f �Ы������t���   ��t�6�Ѓ��    ^]����������������U��h@��uh�f 苫����]�������U��E�D�� ]��U��EHV����   �$� S�   ^]áT�@�T�����   �u������=�6  }�����^]Ëu��t�jh0�jmj�+H������tl����J���P���tfV���\O���   ^]��u�u�9����������H^]�^]�t����T�u.����������5P���t���aK��V�[H�����P�    �   ^]Ã��^]�0R�R�R(R�R�R��������U���Mu�E�H��E�L��   ]� ���������������U��hX�jh�f ��������t
�@��t]�����]�������U��VhX�jh�f ����������t=�~ t7�u8�E�u4�u0�u,�u(����P�?J���u�F�Ѓ�4�M���jJ����^]ÍM����ZJ����^]������U��hX�jh�f �|�������t
�@��t]��3�]��������U��hX�jh�f �L�������t
�@��t]��3�]��������U��hX��uh�f ������]�������U����p�V���.�vf(�fTP�f(�f/�fTP��U��M��M��  f/��  ���f/�vFf/�v@�,��,���   ��$    ������ʅ�u�fn�����^��^��.�v^��]�f/�v(��(�����^��%��f/�v1(��Y��Y��Y��.�E�(��Y��v(��M��M�f/�v(��f�E��E���    �E��E��O+  �M��]��E�f/��f��M��E��E�s�f^�^��]�W������F^��]����U���E���f/�V��w���f/�v(��Y�����X���E�E�$�G  ��������F�������^]� ���U����M3��UW�f/�V��fTP��X����3�f/��M��E���3�;������M�$�+G  �EfTP��E�X����E�E�$��F  ������]�Ef/��Fv'�D�hx�j�@��0  ��������F�} u�fW`�����-�����^��]� ����U���E���f/�V���Fv'�D�hx�j,�@��0  ��������F^]� ������U���M�����f/�V��v'�D�hx�j5�@��0  ��������M����Y��E��E��$��E  �]��F�$��E  �E��]��^E��E��E��$�E  ��E�$�E  �����^�-���^��]� �����̡D�Q�@D�@$�Ѓ����������������U��D�j �u�@D� �Ѓ�]��������U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@D�@�Ѓ���������������̡D�Q�@D�@�Ѓ���������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ����������������U��D��@D� ]��U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ���������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ����������������U��D��uh2  �@D� �Ѓ�]�����U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ���������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ���������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ���������������̡D�Q�@D�@�Ѓ����������������U��D�j �u�@D� �Ѓ�]��������U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ����������������U��D��uh'  �@D� �Ѓ�]�����U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ����������������U��D��uhO  �@D� �Ѓ�]�����U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��D����@XQ�M�Q� �ЋM���o ��~@��f�A��]� ���������U��D����@XQ�M�Q�@�ЋM���o ��~@��f�A��]� ��������U��D����@XQ�M�Q�@�ЋM���o ��~@��f�A��]� ��������U��D���`�@XQ�M�Q�@�ЋM���o ��o@�A�o@ �A �o@0�A0�o@@�A@�o@P���AP��]� U��D��uQ�@X�@�Ѓ�]� �����U��D��uQ�@X�@�Ѓ�]� �����U��D��uQ�@X�@�Ѓ�]� �����U��D��uQ�@X�@�Ѓ�]� �����U��D��uQ�@X�@$�Ѓ�]� �����U��D��uQ�@X�@ �Ѓ�]� ����̡D�j h�  �@D� �Ѓ�����������U��D�V�u�@@�6�@�Ѓ��    ^]��������������̡D�Q�@D�@(�Ѓ���������������̡D�Q�@D�@�Ѓ����������������U��D��u�u�@DQ�@�Ѓ�]� �̡D�j h:  �@D� �Ѓ�����������U��D�V�u�@@�6�@�Ѓ��    ^]���������������U����D��U��E�    �E�    R���   j�@�����#E���]�����������̡D�j h�F �@D� �Ѓ�����������U��D�V�u�@@�6�@�Ѓ��    ^]���������������U��E����u��]� �E��U��D��E�    Rj���   �@������؋�]� ̡D�j h�_ �@D� �Ѓ�����������U��D�V�u�@@�6�@�Ѓ��    ^]����������������    ���A    �A    �A    ���V��V��:���FP��:�����F    �F    ^������������U��V��W�}j�    �F    �F    �F    �G;Gu2j�   ��tY�����G�A��G_�A�F�    ��^]� j�   ��t'�����G�A��G�A��G�A�F�    _��^]� �����U��V�u���    �F    �F    �F    �  ��^]� U��V�u���  ��^]� �����������U��SV��V��9���FP��9���]���F    �F    ��t(�D�h��jI�H��    P���   �Ѓ����u^3�[]� W�}��t;�D�h��jN�H��    P���   �Ѓ��F��uV�K9����3�_^[]� �~�   _�^^[]� �������������V��V�9���FP�9�����F    �F    ^������������U��SV��WV��8���^S��8���}���F    �F    ����   �? ��   �W����   �D�h��jl�H��    P���  �Ѓ����t<� t?�W��t8�D�h��jq�H��    P���  �Ѓ����u���%���_^3�[]� �G�F�G�F��P�7�6�s;  �����t�F��P�wQ�Z;  ��_^�   []� �����������U��SV��WV��7���~W��7�����F    �} �F    ��   �]����   �D���    h��h�   Q�@���  �Ѓ����t?�} tJ�U��tC�D�h��h�   �H��    P���  �Ѓ����u���)���_^3�[]� �E�F�,�F   �D�h��h�   j�@���  �Ѓ����t���    �^P�u�6�G:  �M����t�F��PQ�7�.:  ���   _^[]� ��_^�   []� ����������������    �A    �A    �A    �����U�������   �U��WɉD$VW�H�L$P�L$H�D$    �<��L$}
��_^��]� �u�}���`  �W�f(�f�$�   ��T$(�@�o$��~\��A(�f��d$X�@�\$@���D��\��|��\ŋD$�\�)l$0�f��L$p����   ��$�   ���D$ �����$�   �D$��	��$    ���\$@�f(��L$x���T$p�@�4��\��d��\��l��\�(��Y��Y��Y��Y�f��\�f(��Y��Y��X\$�\��od$X�\��\$�X|$ �t$p�XT$((�f�(l$0�L$ �T$(J�S������$�   ��$�   �L$ �\$W��f�F(��Y�(��Y��X�f(��Y��X��4  �L$W��T$ �|$(f.ş��Dz	W�f(��2����^�f(��Y��D$pf(��Y��Y��D$xfD$p�FHf�^X�P�fT�fT�f/���   f(�fT�f/���   �FH�VX(��fP(��Y��Y��Y��\��\��\�f��^f�f(�~P�NX(��n (��YV(�vH�Y��\�(��YF(�Y��T$0�Vf(��Y��Y��\��   fT�f/��VX��   �FP�NH(��Y��Y��\��\��Y��\�f��^f�N(�f(�n (��YNP(��YFX�vH�\�(��Y��Y��L$0�Nf(��YNP�Y^X�\��\��oD$0f��F0f�v@�   �NPf(��Y�(��Y��\��FH�Y����\��\�f��^0f�F@(��fX�YF@(��YN8�v0�\�(��Y��Y��L$0�NHf(��YN8�Y^@�\��\��oD$0f��Ff�v(��$�   VP��.���U���o ��o@�F�o@ �F �o@0�F0�o@@�F@�o@P�D$�FP3Ʌ�~w��rr�@�D$��%  �yH���@�T$W�)D$foʋD$���$    ��o�f���oD���f��;L$|�f��fo�fs�f��fo�fs�f��f~L$�D$     �D$    ;�}s��+���|A�D$�@�D$�B��t$�D$ 3�3����$    �|���;L$ |��u�|$�}�D$ ;�}�D$�T$�@��T$�U�D$ D$�L$���L$�D$�F0�V �D$@� �D$�~(�v@(ϋ��@�YD����d�f(��Yn�Y��Y��X.�XV�XN�X��FH�Y��X��F8�YD��X��FP�Y��X�(��YD��D$f�D��X��FX�Yč@�$��\��X��T�(ËD$�l$X�n0f�L$h(��YN�@�Y��X��3��T$�D$ �X�(��YFH�X�(��YF8�Y��L$0(��Y��YN �o|$0�Xf�XN�X��X�(��YFP�YVX�X��X�f�f�d$(���  ���f(��|$�D$ы��@���T�f(��Yv(��\��YŋD$ �X6�n @�Y�D$ �Y�(��X�(��YFH�Xn�Xff��X��F8�Y��X��FP�Y��X��F@�Y��T$`�X��FX�Y�(��\��\��X�f(��\��Y��Y��YD$X�|$X���X�f��l$@�X��X\$P(��D$P�D$H�~D$(f�D$hf�d$(;D$������D$H_^��]� ���U�������������U�   @t������@��wg�$�n�E� ����E� ���]� �E�
��E�J�]� �E�J��E�J�]� �E�J��E�J�]� �E�J��E�
�]� ���m�m�m�mn����U��S��VW�����%�����   @t�����ʃ��};�t�����t�u�����t��u;�t?�����t7�΁����Eǃ��t����   �_�^�[]� ��   ���Ё�   @�_^[]� �U������4�AW��$W��T$SfD$ V�\$,�L$$�\$�L$W���S  �9�u��$    ������Ш�)  ���������U��Z�@�[�<��l��\<��\l�;Zuc�\��B�\\��@�d��\d��T��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��Xd$(��d�d��B�\d��@�B�@�T��\��\\��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��X\$�XL$�Y��Y��\$�L$�\��Xt$ (��T$ ���L$�����f(��Y�f(��Y��X�f(��Y��X��D+  f(�W�f.П��D�Ez �@_^[��]� ����^�_^[(��YD$� (��YD$�@�D$�Y��@��]� U���<(@��A�=���%8�V�E�3��E�(p��E܅��  �m��u��U��E�S��MW��    ������Ш�n  ���������U��@��tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��EċB�@��tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��Eċz���tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��EċB;���   �@��tU��f/�vf(��\�f/�vf(��\�f/�vf(�f/�vf(��L�f/�vf(�f/�v=f(��7�o��   �~d��E��o��m�f��u��E��U��Eă��M��u���_[��ta�Ef(�f(��X�����X�f(��X�^�Y��Y��Y�f��f�P�\0�\h�\`�Ef��0f�`��]� �EW�W�^� f�H�E� f�H��]� ��������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}���x(���t"�v3Ʌ�~�I ���%���;�tA��;�|�_���^]� _��^]� ���������U��SV�q2�3҅�~9W�9����%���;Eu ����   @u�����t	�   ���3�
�B;�|�_��^��[]� ������������V�q3҅�~�	�d$ ��   @u	�����tB��Nu��^�����V�q3҅�~�	�d$ ����ШtB��Nu��^�����������U���V��3�9N~��$����A;N|�N��~kS�   3�W�U��]�����x:�������;�}+�I ����<����������;�u��   ��@;F|ۋU��]�B�N���]��U��B�;�|�_[^��]�����������h\�jh_� ��������uË@����U��V�u�> t/h\�jh_� �Æ������t��M�M�@Q�Ѓ��    ^]���U��Vh\�jh_� ��艆������t�@��t�u����^]� 3�^]� ��������U��Vh\�jh_� ���I�������t�@��t�u����^]� 3�^]� ��������U��Vh\�jh_� ���	�������t�@��t�u���u�u��^]� 3�^]� ��U��Vh\�jh_� ���Ʌ������t�@��t�u����^]� 3�^]� ��������U��Vh\�j h_� ��艅������t�@ ��t�u����^]� 3�^]� ��������U��Vh\�j$h_� ���I�������t�@$��t�u����^]� 2�^]� ��������Vh\�j(h_� ����������t�@(��t��^��3�^������Vh\�j,h_� ���܄������t�@,��t��^��3�^������U��Vh\�j0h_� ��詄������t�@0��t�u����^]� 3�^]� ��������U��Vh\�j4h_� ���i�������t�@4��t�u���u��^]� ���^]� ����Vh\�j8h_� ���,�������t�@8��t��^��3�^������U��Vh\�j<h_� �����������t�@<��t�u����^]� ���������������U��Vh\�j@h_� ��蹃������t�@@��t�u����^]� ���������������U��Vh\�jDh_� ���y�������t�@D��t�u����^]� 3�^]� ��������U��Vh\�jHh_� ���9�������t�@H��t�u����^]� ���������������Vh\�jLh_� �����������t�@L��t��^��3�^������Vh\�jPh_� ���̂������t�@P��t��^��3�^������Vh\�jTh_� ��蜂������t�@T��t��^��^��������Vh\�jXh_� ���l�������t�@X��t��^��^��������Vh\�j\h_� ���<�������t�@\��t��^��^��������U��Vh\�j`h_� ���	�������t�@`��t�u���u��^]� 3�^]� �����U��Vh\�jdh_� ���Ɂ������t�@d��t�u���u��^]� 3�^]� �����U��Vh\�jhh_� ��艁������t�@h��t�u���u�u�u�u��^]� ���U��Vh\�jlh_� ���I�������t�@l��t�u���u�u��^]� 3�^]� ��U��Vh\�jph_� ���	�������t�@p��t�u���u��^]� 3�^]� �����U��Vh\�jth_� ���ɀ������t�@t��t�u���u��^]� 3�^]� �����U��Vh\�jxh_� ��艀������t�@x��t�u���u��^]� 3�^]� �����U��Vh\�j|h_� ���I�������t�@|��t�u����^]� 3�^]� ��������U��Vh\�h�   h_� ����������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh\�h�   h_� ���������t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh\�h�   h_� ���f������t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh\�h�   h_� ���������t���   ��t�u���u�u�u��^]� 3�^]� ���������U��Vh\�h�   h_� ����~������t���   ��t�u����^]� 3�^]� ��U��Vh\�h�   h_� ���~������t���   ��t�u����^]� ���������U��Vh\�h�   h_� ���F~������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh\�h�   h_� ����}������t���   ��t�u���u�u��^]� 3�^]� ������������U����M�U�E�A�R�X�\B�\��\Y�Y �Y�Y�X��X��U��E���]�����U��h\��uh_� �[}����]��5p�����t��jj �{9  YY�9  U��� SW3ۍ}�j3��]�Y�9Eu��I  �    �;  ����M�E��t�V�E�E��EPS�u�E��E����P�E�B   ��<  �����M�x�M����E�PS�;  YY��^_[��]�;�u����I  ̺0��aK  �0���J  ���������z�����������������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̃��\$�D$%�  =�  ��  �<$f�$f��f����  f$f%Pf`fW�fX��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU�fV�f($������X��\��Y��Y��Y����X��^�ff-��\�fs�?��fs�?�Y�fp�Df5 �Y��Y�fW��Y�f\%��Y��X��Y��\�fp���X��\��\ă��-�  ��A�   fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<���Y��Y��Y��\�fT��X��\��X�f-��\��X�f�^�f fXՐ����Y��Y��Y��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fWƃ���;  = 8  ��   f�f(5f�f( f(%0fY�f(-�fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��XŃ��-�;  ����   fW�fT=Pf%hf(�Y�f( �\�f(0fp�D�Q�fY�fp�Df��fY�fX�f�fY�����Y�fX�fp�D�Y�fT�fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^�fX�fY�fp���X�% �  f��fp���X��X��X��X�fWƃ���� = � ��   f~�fs� f~�������  �?+���� ttf$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�1K  fD$�� �f������fn�fp� f�f�fT�fT��X��f�f��X��fW��Xƺ�  �t���f�$�<N  �$�~$��Ð���\$�D$%�  =�  ��  �<$f�$f��f����  f$f�f(�fT�f/��p  �8  f/�sgf/���  f(�fY�f(�fY�f(-�fY�fX-pfY�fX-`fY�fX-P�Y�f(�f���X��Y��\Ń��f/���   f(�fY�f(�fY�f(-@fY�fX-0fY�fX- fY�fX-fY�fX- fY�fX-�fY�fX-�fY�fX-��Y�f(�f���X��Y��\Ń���~�fW�f/�sO�~��~-��~��X�fs�,f��f~؍@�~,�ȅ�~��\��Y��X��^�f���   �~��~��^�f��~Ÿ��~$���f(�fY�f(�fY�f(-�fY�fX-pfY�fX-`fY�fX-P�Y�f(�f���X��Y��\��\��\�fVƃ��f/�u	f$���f/�sf$�Y҃��f$f��Y҃���~��~�fT�f.�z�D$��f��X����ú�  ���T$�ԃ��T$�T$�$��G  fD$���f�$�L  �$�~$��ÍI �������̃��\$�D$%�  =�  u�<$f�$f��f���d$�n  f��f%�f-00f=��6  f0�Y�f8�-��X�fP�\�f(@�Y�fɁ�v ����?f(- �����fY��\��YX�\�fxf����\�fY�f\�f(5 �Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�Y fX5�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��f��f%�f��f��\�f(�Ã�f�$��K  �$�~$����������̃��\$�D$%�  =�  ��  �<$f�$f��f����  f$f�f( f(5�f(f( f��%�  ��@  +�-�<  Ё�   ��  fY�fX�f(�f\�fY�f(%0fY�f(-@f\�f~��ȃ�?������f\�f(�PfY�f(�fY�fX��Y��X�f�fo5�f��fo5�f��fs�.fY��X�fV�f��X���~  ��|  w�Y��X�Ã���|$f�T$f�� f�$�,$����+�fo5�f���  fn�fs�4fV���  fn�fs�4f$�$ft$�D$����f$$�$���$f$�l$��f�����  ���  s*�� t,��Á�   �r��+#��wr�$���9��s��ú   ��   ��fD$�T$�ԃ��T$���T$�$��C  fD$�� �=  �s1�D$=   �sf� �Y��   �f� �Y��   뙋$=  �w(�� u#�D$=  �ufp ���fx ��ú�  �]����D$%���=  �@�x���f$�XP ���f�$�#J  �$�~$��Ã��\$�D$%�  =�  �8  �<$f�$f��f���#  f$fL$f=0Yf@YfT���fs�,f�� fV�f��%�   ��%�  �Y<�� f,�� �f(4��$��  +у�ʁ�   ���  �    �� fn�f��fs����f�Y��fs�&f�� fT%0Y%�   ��%�  �Y��,�Y,��,�fX4��0fV%@Y�X�fT���fs�f�� f�Y�\�f=�Y%�  ��%�  �Y,��8�Y��8fX4��@fT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�f�Yf���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%�YfT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f( Q�Y��-��Y�f(Q�X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X YfY��\ YfY��\�����f(� Qf(5`YfY�fX�fp���Y�fW���?  �X�f���X�f%�Yfn��YT$�Y�fs�-fp�Df(=pY�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��X��X��X��XÃ��fL$fPYf~���fT�fs� f~Ɂ�  ���   ��� �B  �� �   �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$f(ѹ�  fn�fTPYfs�4f��f�Yf��fv�f��%�   �� ȁ�   ��r[�� f0Yf@Y�5���f<$f(�f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=0Yf@Y�Y�f~�fs� f~��� tRfT���fTPYfs�,f�� fV�%�   ��%�  �Y<�� f,�� �f(4��$�> �n����Ё������ u��T$��   ��� t0��#��  ��fn�fs� f@Yf$�^ʺ   �  ��#��� ��   fW����f0YfW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   umfL$f(ѹ�  fn�fTPYfs�4f��f��f��fv�f��%�   =�   t-fL$f��% �  �� tf�Y���f�Y���fL$f��% �  �� �a  fW����fL$f��% �  �� �@  fW�����X��ĺ�  �  f$f~�fs� f~ҁ����¹    �� �k���f�Yf�Y�Yɺ   �Q  f$$fT$f0YfW�fT�fv�f��%�   =�   ��   f~��� u)fs� f~��  �?��   ��  �uf@Y���f0YfW�fT�fv�f��%�   =�   ucf��f$$% �  ��  �у� ��   �� tf��%�  =�?  r!fW����f��%�  =�?  sfW����f�Y����X��º�  �Vf~�fs� f~��������f@Y�   �� t-f~�   %���=  �wr�� w���f� �   ��fD$�T$�ԃ��T$���T$���$�:  fD$��(Ã� ~(=   �"  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X Y���� fY��\ YfY��\�����f(� Qf(5`YfY�fX�fp���Y��X��X�f%�Yfnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(=pY�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� A^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� � ������^�X��Y��Y��X�f��%�  �   =�  ������   �� ��������f�Yfn��Y�fs�-fV��   �����   �� tf�Y�Y�Y�}���f�Y�Y��l���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r�ɀ� fn�fs�-���f$$f�����  ���?  f��3�% �  �� �;����Y���f�$f�L$�`?  �$�~$��Ã��\$�D$%�  =�  u�<$f�$f��f���d$�{  f��f%�f-00f=��6  f b�Y�f(b�-��X�f@b�\�f(0b�Y�fɁ� v ����?f(-b��Y���fY��\��YHb�\�fxf����\�fY�f\�f(5�a�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX- b�Y fX5�afY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��,f��f=�u	�Y`b�fPb�Y��\��YXbÃ�f�$�&@  �$�~$��ÍI �������̃��\$�D$%�  =�  ��   �<$�$������   f����%�  =�  t0��% �  u�Q����f�$�<$ uP�� �  uHf���� u>�ً���u$f��%��  uf��%��  uf�� %��  t�f�$�L$��  ��$    �D$  ���1   ���T$�ԃ��T$�T$�$��4  fD$���f�$��?  �$�~$��Ë��=�� �l@  ���\$�D$%�  =�  u�<$f�$f��f���d$�;@  � �~D$f(�bf(�f(�fs�4f~�fT�bf��f�ʩ   tL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�4  ���D$��~D$f��f(�f��=�  |%=2  �fT�b�X�f�L$�D$���b�f��bfT�bf�\$�D$���̃=�� �#@  ���\$�D$%�  =�  u�<$f�$f��f���d$��?  � �~D$f(�bf(�f(�fs�4f~�fTcf��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$��2  ���D$��~D$f��f(�f��=�  |!=2  �fT�b�\�f�L$�D$����f� cfV cfT�bf�\$�D$����������������WV�t$�L$�|$�����;�v;��h  �%��s��  ���   ��  ��3Ʃ   u�%����  �%�� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����H�����   u������r*��$�H���Ǻ   ��r����$�\��$�X���$�ܡ�l�����#ъ��F�G�F���G������r���$�H��I #ъ��F���G������r���$�H��#ъ���������r���$�H��I ?�,�$��������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�H���X�`�l����D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�������$����I �Ǻ   ��r��+��$���$������D��F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ������������ȣۣ�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������� ��D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋T$�L$��t�D$�%��s�L$W�|$��]�T$���   |�%���E9  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�Q�$c�@:  Y�U��V��������EtV�K���Y��^]� U���   �} t�E  ��]ø����������*������ �	��$��(����,�B��0����4����jh@���Y  �E��uz�M  ��u3��F  ��H  ��u�|M  ���GY  �����T  �h��cM  ��y�5I  ���YP  ��x �R  ��xj �J  Y��u�d���   ��O  �Ʌ�ue�d���~�H�d��e� �=�� u�nJ  �@I  �u��u�O  ��H  ��L  �E������   �   �u��u�=8��t�H  ��p��u^�58��+T  Y��u[h�  j�W  YY���������V�58��!T  YY��tj V�*G  YY����N��V�t  Y�������uj �EF  Y3�@�X  � U��}u�LR  �u�u�u�   ��]� jh`��+X  3�@�u��u95d���   �e� ��t��u5�,c��t�uV�u�щE����   �uV�u�����E����   �]SV�u腪�����}��u(��u$SP�u�m���SW�u������,c��tSW�u�Ѕ�t��u*SV�u�������#��}�t�,c��tSV�u�Ћ��}��E��������&�M�Q�0�u�u�u�   ��Ëe��E�����3��oW  �U��}u�uj �u�G����u�u�C  YY]�U��} t-�uj �5������uV�   ����P��   Y�^]�U��V�u���woSW�����u��X  j�-Y  h�   �F  ���YY��t���3�AQj P������u&j[9(�tV�`X  Y��u���>   ��7   ���_[�V�?X  Y�#   �    3�^]�����������WV�t$�L$�|$�����;�v;��h  �%��s��  ���   ��  ��3Ʃ   u�%����  �%�� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����h�����   u������r*��$�h���Ǻ   ��r����$�|��$�x���$��������ܬ#ъ��F�G�F���G������r���$�h��I #ъ��F���G������r���$�h��#ъ���������r���$�h��I _�L�D�<�4�,�$���D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�h���x��������D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�������$����I �Ǻ   ��r��+��$���$����<�d��F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ����ȮЮخ�����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$������,�@��D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̺���  ���<  �����������̃��\$�D$%�  =�  �  �<$f�$f��f����  f$f%�zf�zfW�f�z��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU@rfV�f($�@c���X��\��Y��Y��Y����X��^�f=�zf-xz�\�fs�?��fs�?�Y�fp�Df5�z�Y��Y�fW��Y��Y��X��Y��X�fp���X��X��Xă��-�  ��C�  �Y��\��Q�f��fs�fT=pzfs���f%�z���\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<�@r�Y�f(@z�Y��Y��\��X��\��X�f-xz�\��X�f�z�^�f�zf\�@c���Y�%�   ���Y��Y��Y��Y��X�f���Y��X�f���X�fp���\��X�fVƃ���;  = 8  s]f�f(5�zf�f(�zf(%�zfY�fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X����-�;  ���B  �Y��\��Q�f��fT=`zfp�DfT`z��f%�z���\��Y��X��Y��\����Y��Y��\��\��X��\�f(�zfp���\��X�fp���X��Y��X�fp���^�f(�zf(-�zf(�zfY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(@z�Y�fX�fp���Y�fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fVŃ���� = � ��   f~�fs� f~�����  �?+���� tpf$f~�fs� f~с��������  ��� }rfW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�@  fD$�� �f�zf@zfHz�X�fU�fV����f$fW��Xƺ�  �f$fW���f�����  �����  r�X�fV��Y����f�$�P  �$�~$��Ë������������̃��\$�D$%�  =�  �Y  �<$f�$f��f���D  f$�    f(�f�fs�4f�� f({f(p{f(% {f(50{fT�fV�fX�f�� %�  f(��{f(� �fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(�{f(�f(�{fY�fY�fX�f(�{�Y�f(-@{fY�f(�P{fT�fX�fX�fY��Y�fX�f(�f�fY�f(�fɃ��X��X��X��f$fW���� f�� �� wL���tb���  wpf$f({f(p{fT�fV���� f�� �� t��f�{ú�  �Ofp{�^�f�{�   �4f�{�Y�������=��������  ���  s<fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$�b  fD$�� �f$f(�f~�fs� f~с��� ��� t���  �f�$��N  �$�~$�������Vjj �F  YY��V� ���������ujX^Ã& 3�^�jh���G  �e� �(:  �e� �u�#   Y���u��E������   ���G  Ëu��:  �U��QSV�5�W�5�����5���E��֋؋E�;���   ��+��O��rvP�O  ���GY;�sG�   ;�s�Ƌ]��;�rPS�sF  YY��u�F;�r>PS�_F  YY��t1��P��� �����u� ��K�Q� �����E�3�_^[��]�U���u�������Y���H]�U��U� ��ҋM#�#Mщ �]��O  ��tj�2O  Y� �t!j���  ��tjY�)jh  @j�   ��j�'8  �U��E�p�]�U���(  ��3ŉE��}�Wt	�u�R  Y������ ������jLj P���������������������0���������������������������������������������f������f������f������f������f������f��������������E�������E������ǅ0���  �@��������E�������E�������E������� ���������P��C  Y��u��u�}�t	�u�"Q  Y�M�3�_������]�U��E�t�]�U���5t�����t]���u�u�u�u�u�   �3�PPPPP��������j��  ��tjY�)Vj� �Vj�s���V�LC  ��^�U��V�uWV�R  Y�N�����u�Y  � 	   �N ����  ��@t�=  � "   ��S3���t�^��t}�F�����N�F���^���F�  u*��P  �� ;�t�P  ��@;�uW�Q  Y��uV�\  Y�F  tz�V�+ʉM�B��FH�F��~QRW��Q  �����G�� �N�h���t���t�ǋ������������@��A tjSSW��Z  #����t%�N�E��3�@P�E�EPW�dQ  ����;]t	�N �����E��[_^]�U��V��M�F ��ufW�H1  ���~�Wl��Oh�N;��t�x��Gpu�^  ��F_;T�t�N�x��Apu�b  �F�N�Ap�u���Ap�F�
���A�F��^]� U���  ��3ŉE��E������SV�������EW�u�}������3��؉������������������������������������������������������������&  ����������������
  �@@ucP�O  Y�ȃ��t���t�������������@��B$��
  ���t���t�������������@��A$��T
  ���������F
  �3��������ȉ���������������������������������	  ������@����������	  �B�<Xw��������3����������(��ǉ����������������������w	  �$���3���������؉������������������������������������<	  �� tF��t9��t/HHt���������	  ���������	  ����������  �����ˀ   ������*u/�������������������  ���؉������������  k�����
�����������  3��������  ��*u+������������������������p  ��������d  k�����
�����������>  ��ItE��ht8��������lt��w�,  ��   �����8lu@��   �������������� ������������ <6u�������4u�ǃ��� �  ����<3u�������2u�ǃ����������<d��  <i��  <o��  <u��  <x��  <X��  3��������3�������������P��P�hb  YY��t8������P�������������  ���������A���������������d  ������P�������������  ����  ��d��  �Q  ��S��   t|��AtHHtVHHtHH�  �� ǅ����   ��������������������@�   ���������������2  ǅ����   �  ��0  ��   ��   �������   ��0  u��   �������������������t�ʋ7����������  �S  ��u�5(�ǅ����   �ƅ�t3�If9t����u�+����<  ��X��  HHtp���'���HH�$  ����������  t0�G�Ph   ������P������P��b  ����tǅ����   ��G�������ǅ����   ��������  �����������t3�p��t,� ��   t�+�ǅ����   ���  3ɉ������}  �5$�V�`  Y�k  ��p��  ��  ��e�Y  ��g�K�����itd��nt%��o�=  ǅ����   ��y[��   �������M�����������`  ���  �������� tf���ǅ����   �z  ��@������ǅ����
   �� �  u��   ��  ���������3����  u��guVǅ����   �J;�~��������=�   ~7��]  W�;  ������������Y��t
���������
ǅ�����   ����������������������G�������������P��������������P������������VP�5(����Ћ�����   t!������ u������PV�54�����YY������gu��u������PV�50�����YY�>-�(�����   F����������ǅ����   j���s�����HH��������k  j'ǅ����   X���������|���Qƅ����0������ǅ����   �^�����3��������� t��@t�G���G����@t
�G���ȋ���O�����@t;�|;�s����߁�   �������� �  u����������y3�B�����   ������;�~�Ћ��u�������u��J�����������t=�������RPWQ�n_  ��0����������������9~������������N������밋������E�+�F��������   t6��t�>0t-N�������0�!��u�5$����I�8 t@��u�+Ɖ����������� ��  ��@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����������+���u������P������Wj �  ��������������������Q������P������P�  ����t��u������P������Wj0�  �������� ������t}��~y��H���������Pj�E􉍄���P������P��]  ����u?9�����t7������������P�������E�������P�t  ����������������u��(����������#������������Q������PV�:  ����������x#��t������P������Wj ��   ����������������tP�����3�Y��������������������������������������������� _^[t
�������ap��M�3�������]��P  �    ���������/�7�k�����c���U��U�B@t�z t/�Jx��M������ER��P�w���YY���u�E��]ËE� ]�U��V�u��~W�}W�uN�u�������?�t���_^]�U��V�uW�}��E�G@t� u
�M�E�N�& S�]��~@�EP�EKW� P�I����E���E�8�u�>*uPWj?�-����E����˃> u�E�[_^]��~$  ��u���Ã��U��V������MQ��    Y���   �0^]��J$  ��u���Ã��U��M3�;�0�t'@��-r�A��wjX]Í�D���jY;��#���]Ë�4�]�U��� �j����A  �u�t4  �=�� YYuj�A  Yh	 ��B4  Y]�U���$  j���  ��tjY�)�x��t��p��l��5h��=d�f���f���f�`�f�\�f�%X�f�-T������E �|��E����E������������  �������x�	 ��|�   ���   jXk� ǀ��   jXk� ���L�jX�� ���L�h���������]�������U���0���S�ٽ\�����=|� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=|� t�#  ��8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����3  �   [�À�8�����=`� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��������������������s4����,ǅr���   ��������������������v���VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�X  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����K   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[��������̀zuf��\���������?�f�?f��^���٭^����܄�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����܄�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����Ԅ���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t���U��%�� ��S3�C	��j
��  ���L  3ɉ��3��V�5��W�}����_�O�W�E�M��E��ineI�E�5ntel�5��ȋE�5Genu���j�X��j Y���_�O�W�M�M�tC�E�%�?�=� t#=` t=p t=P t=` t=p u�=�����=����=���}�|5j3ɍu�X���Ƌ5���X�H�M��P�E�   t���=���3���   tM�����   �5����   t2��   t*�����   �5��� t�� ���   �5��_^3�[��]�U���(3��E��E�9��t�5 ����������E��   V;���  ��  ���  ��   jZ+���   H��   ����   H��   ����   HtN��	�#  �E�   �E�h��E�u� �E�]�� �E��]��P�]���Y����  ������ "   ��  �E�d��E�u�E�   � �E�]�� �E��]��P�]���Y�  �E�   �E�d���E�\��V  �U��E�\��l����E�X��;  �U��E�X��Q����E�h�놃�tfHtWHtHHt/���  ��	t���8  �E�l���   �E�t���   �E�h��E�u� ���   �E�h���   �E�   ������E�����   �E�   �E�|������������   �$�C��E�X���E�\���E�d���E܄���E܌��u����Eܔ��i����Eܜ��]����Eܤ��E�u� �M��� �E�]�� �]��.�Eܨ����Eܬ����Eܰ��E�u� �E�]�� �]���E��E�   P�]���Y��u����� !   �E��^��]À�����������4�����������������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��R  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�R  ���$��X  �   ��ÍT$�mX  R��<$tmf�<$t�)X  =  �?s-����������������=`� ��X  �   ����X  w8�D$��%�� D$u'��   ���t���������W  ���� u�|$ u����-���   �=`� �*X  �   ����3W  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��X  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�X  ���$�rW  �   ��ÍT$�W  R��<$t6f�<$t�-������=`� �PW  �   ����MW  ��V  �&��� u�|$ u����-ʄ�   �t���뻸   �=`� �W  �   ����V  Z������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�Z  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�UZ  ���$�RV  �   ��ÍT$��U  R��<$tPf�<$t�-��������z�=`� �,V  �   �б�)V  �-����������z��������U  ���� u�|$ u����-���   �=`� ��U  �   �б��T  Z�������̃=�� tn���\$�D$%�  =�  u�<$f�$f��f���d$uA�-[  ��=�� t<���\$�D$%�  =�  u�<$f�$f��f���d$u��Z  �Z��9����Z��c�������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uZ�Z_  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�_  �����$�T$�D$�   ��ÍT$�8T  ��P��<$f�<$t��S  ��  ��T$��  ���   �	T  ��   �  ���   �L$���S  ���S  ��u���=`� �)T  ���   �dT  �=`� �T  ���   ��R  ZÍT$�S  �D$uA�3���   ���D$u����   �3��3�%�� D$uÍT$�[S  �D$��%  ����� =  �uT$u���u���t��Q���$�\$��q�i  ��Y�a���t���eS  �   �B����D$%�� D$������؋D$%���D$t=�f   �l$���D$�   t�- ���t��   ���������S  ����R  ������R  ���   ��������������-���   ���������ٱ ����u���������ٛ���u�����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��i  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�ui  ���$�R  �   ��ÍT$�Q  R��<$tPf�<$t�-��������z�=`� ��Q  �   ����Q  �-����������z��������?Q  ���� u�|$ u����-���   �=`� ��Q  �   ���P  Z�������̃��$�MQ  �   ��ÍT$��P  R��<$�D$tQf�<$t�P  �   �u���=`� �#Q  �   � �� Q  �  �u,��� u%�|$ u���P  �"��� u�|$ u�%   �t����-���   �=`� ��P  �   � ���O  Z�j
��  ���3��U��QQSV���  V�5��r  �E��YY�M��  ��#�QQ�$f;�uT�q  YY��~-��~��u#�ESQQ�$j�Pl  ���qVS�Jr  �EYY�c�E���S�����\$�$jj�?�0i  �U��E��������DzV��S���r  �E�YY��� u�S�����\$�$jj�7i  ��^[��]�U��QQSV���  V�5���q  �E��YY�M��  ��#�QQ�$f;�uT�p  YY��~-��~��u#�ESQQ�$j�yk  ���qVS�sq  �EYY�c�E���S�����\$�$jj�?�Yh  �U��E��������DzV��S���.q  �E�YY��� u�S�����\$�$jj�`h  ��^[��]Å�uf���fn�f`�fa�fp� SQ�ك���ux�ڃ���t0ffAfA fA0fA@fAPfA`fAp���   KuЅ�t7����t��I f�IKu���t����t
f~�IJu���t�AKu�X[��ۃ�+�R�Ӄ�t�AJu���t
f~�IKu�Z�^���̋T$�L$��   u@�:u2��t&:au)��t��:Au��t:au������uҋ�3���������Ë���   t���:u����t���   t�f���:u΄�t�:auń�t����jh���   j�p  Y�e� �u�F��t0�������M��t9u,�A�BQ�����Y�v�����Y�f �E������
   �   Ë���j�q  Y�U��j �u�u�u�u�u�u�   ��]�U��E��et_��EtZ��fu�u �u�u�u�u��  ��]Ã�at��At�u �u�u�u�u�u�}  �0�u �u�u�u�u�u�   ��u �u�u�u�u�u��  ��]�U���,SVWj0X�u���E��  �M�3ۍM������}��y���u��t�M��u	����j��G�;�w����j"_�8�������  �U��Z�E����%�  =�  uy3�;�uu���;�t�A�j WP�^SR��  ������t� �  �;-u�-F�}��j0X�����$�x�F�FjeP�us  YY��t�����ɀ����p��@ 3��O  3���   ��t�-F�} �]j0X�����$�x�ۈF�Jۃ����  ���'3���]�u'j0X�F���B�
%�� �u3��E���E��  ��F1����F�M��u� ��Eԋ��   � � ��B%�� �E�w	�: ��   �e �   �E��M��~S��R#E#ыM����� ����w  j0Yf�����9vËM�U�F�E���E�E�����O�M�E�f��y�f��xW��R#E#ыM����� ���w  f��v6j0�F�[���ft��Fu�H��]�;E�t���9u��:��	�����@���~Wj0XPV��������E�8 u���} �4�U����$�p���R�!w  �ȋ�3����  #�+M��x;�r	�F+����F-��������0��;�|A��  ;�rPRSQ��u  0�U�F3�;�u;�|��drPjdSQ��u  0�U�F3�;�u;�|��
rPj
SQ�u  0�U�F�]�3���0����F�}� t�M܃ap���_^[��]�U��j �u�u�u�u�u�V  ��]�U����M�SW�u �5����]��t�} w	�K���j��U3����ǃ�	9Ew�-���j"_�8�q�����   �} t �M3�����P3��9-���P��  �UYY�EV��8-u�-�s��~�F�F�E����   � � �3�8E�������9Et��+�EhȝPV��j  ����uv�N9}t�E�U�B�80t-�RJy���F-jd[;�|��� Fj
[;�|��� F V���^t�90uj�APQ�4������}� t�M��ap���_[��]�WWWWW�~����U���,��3ŉE��E�M�S�]VW�}j^VQ�M�Q�p�0�Hs  ����u������0�(������t�u��u
�����j^����;�t3��΃}�-��+�3�����+ȍE�P�CPQ3Ƀ}�-��3�������P�p  ����t� ��u�E�j P�uSVW��������M�_^3�[������]�U����E�M�SV�u�@H�E������u��t�} w�"���j[��f����   3�W�}8]t�M�;�u�U3��:-���f�00 �E�8-u�-F�@��jV�  Y�0FY����~JjV�  �E�YY���   � � �F�E�@��y&8]t�������;�|��WV�l  Wj0V蠽����_�}� t�M�ap�^��[��]�U���,��3ŉE��E�M�SW�}j[SQ�M�Q�p�0�q  ����u�+�����r������lV�u��u������Z������S���;�t3��΃}�-��+ȋ]�E�P�E��P3��}�-Q���P�nn  ����t� ��u�E�j PSVW�g�����^�M�_3�[�:�����]�U���0��3ŉE��E�M�SW�}j[SQ�M�Q�p�0��p  ����u�j�����������   V�u��u�O�����������   �E�3�H�}�-�E�������9;�t��+��M�Q�uPS�m  ����t� �S�E�H9E������|+;E}&��t
�C��u��C��u�E�jP�uVW��������u�E�jP�u�uVW�I�����^�M�_3�[�;�����]�U��j �u�   YY]�U���W�u�M��Z����U�}��
��t���   � � :�tB�
��u��B��t4�	<et<EtB���u�V��J�:0t����   ��:uJ�BF���u�^�}� _t�E��`p���]�U��j �u�u�u�   ��]�U��QQ�} �u�ut�E�P��m  �M�E���E��A��EP�Dn  �M�E�����]�U��j �u�   YY]�U����M�V�u�o����u�P�j  ��e�F�P�Bi  ��Yu��P�j  Y��xu���E�����   � � �F���ȊF��u�^8E�t�E��`p���]�U��E�������Az3�@]�3�]�U��W�}��tV�uV��8  @P�>VP������^_]�Vh   h   3�V��o  ����u^�VVVVV�+����V3����� ��������(r�^�U��V��  �����E  �V\��W�}99t�����   ;�r�   ;�s99t3Ʌ��  �Q���  ��u�a 3�@��   ��u�����   �ES�^`�F`�y��   j$_�F\�d �����   |�9�  ��~du�Fd�   �   �9�  �u	�Fd�   �u�9�  �u	�Fd�   �d�9�  �u	�Fd�   �S�9�  �u	�Fd�   �B�9�  �u	�Fd�   �1�9�  �u	�Fd�   � �9� �u	�Fd�   ��9� �u�Fd�   �vdj��Y�~d�	�q�a ��Y�^`���[�3�_^]�U��csm�9Eu�uP����YY]�3�]�jh���J  �u����   �~$ t	�v$�-���Y�~, t	�v,����Y�~4 t	�v4����Y�~< t	�v<� ���Y�~@ t	�v@����Y�~D t	�vD����Y�~H t	�vH�ӻ��Y�~\Нt	�v\�����Yj�/c  Y�e� �Nh��t�����u��0�tQ薻��Y�E������W   j��b  Y�E�   �~l��t#W�e-  Y;=��t����t�? uW��+  Y�E������   V�>���Y�  � �uj�d  YËuj��c  Y�U��8����t'V�u��uP�l  ��8�Yj P�{  YYV����^]�V�   ����uj�  Y��^�VW���58����$  ��Y��uGh�  j�  ��YY��t3V�58��  YY��tj V�%   YY���N���	V�o���Y3�W�$�_��^�jh��X  �u�F\Н�f 3�G�~�~pjCXf���   f���  �Fh0����   j�a  Y�e� �Fh�����E������>   j�la  Y�}��E�Fl��u����Fl�vl��)  Y�E������   �  �3�G�uj�b  Y�j�b  Y��  �Jb  ��u�c   3��h
��  �8�Y���t�Vh�  j�R  ��YY��t-V�58���  YY��tj V�����YY���N��3�@^��   3�^á8����tP�r  �8��Y��`  U��Q�E�Php�j �,���th���u��0���t�u�Ћ�]�U���u�����Y�u�(��VW�5�����5������t�> t�6誸��Y��u�5��SV藸���5��3ۉ��Y��t9t�6�y���Y��u�5��V�g����5������V����5���K��������������;�t9��tW�'���YV� ����� ���tP����Y� �����tP�����Y���T���0N[u�T��0�;�tP�ͷ��Y�5T�_^�U����  �u�;  Yh�   �   �jj j �>  ���U��=(c th(c�j  Y��t
�u�(cY����h�h���   YY��uCh4 �����$ �h���v   �=�� YYth���i  Y��tj jj ���3�]�U��j j�u�   ��]�Vj � ���V�  V�����V����V�  V�j  V�j  ��^��	  U��ESV�u3�+ƃ���9uW���#�v���t�Ѓ�C;�r�_^[]�U��V�u3����u���t�у�;ur�^]�j��]  Y�j�@_  Y�jh��V  j��]  Y�e� �=����   ���   �E����} ��   �5���5��֋؉]ԅ�tt�5���֋��]�}��}܃��}�;�rWj � �9t�;�rG�7�֋�j � �����5���5��։E��5���֋M�9M�u9E�t��M�ى]ԉE����h0�h �����YYh8�h4�����YY�E������    �} u)���   j�-^  Y�u�^����} tj�^  Y��y  ��<�3ɣ��������Ã%�� �jdh0��
  j�u\  Y3ۉ]�j@j _W��
  YY�ȉM܅�uj��E�Ph���]  ������[  ����=��   ;�s1f�A 
�	��Y�a$��A$$�A$f�A%

�Y8�Y4��@�Mܡ���ƍE�P�L�f�}� �/  �E����$  ��M���E���E�   ;�|�ȉM�3�F�u�9��} j@W�
  YY�ȉM܅���   ����M���}�j�[�E؋U�;���   �2���t[;�tW� �tQ�uV�D��U���t<����������4����u܋��E؊ �Fj h�  �FP�V  ���F�U��M�G�}ԋE�@�E؃��U�냉���=������   ;�s$f�A 
�	��Y�a$�f�A%

�Y8�Y4��@�M���F�uЋM�� ���j�[3��}ԃ���   ����5���u܃>�t9t�F��F�   �F���uj�X�
�G�������P�@��E���tL��tHP�D���t=�M�%�   ��u�F@���u	�F�Fj h�  �FP�J  ���F��F@�F��@���t���XG�=����]��   3��	  �j�@[  Y�VW����>��t7��   ;�s"���� tW�H����@��   �G�;�r��6�����& Y������|�_^�U��QQ�=�� u�\%  SVWh  ���3�WS����P��5��=����t8u���E�P�E�PSSV�]   �]��������?sE�M����s=��;�r6R�  ��Y��t)�E�P�E�P��PWV�    �E���H�=�����3�����_^[��]�U��ES�]V�uW�# �}�    �E��t�8���E3ɉM�>"u3�����F�Ȱ"�M�5���t��G�F�E��P�+e  Y��t���t��GF�E��t�M��u�< t<	u���t�G� �N�e �> ��   �< t<	uF��> ��   �U��t�:���U�E� 3�B3��FA�>\t��>"u3��u�} t�F�8"u���3�3�9E���E���I��t�\G���u���tA9Mu< t8<	t4��t*��P�Xd  Y��t��t��GF���G���tF��F�o�����t� G��-����U_^[��t�" �E� ]Ã=�� u�2#  V�5h�W3���u����   <=tGV�R*  FY����u�GjP�v  ���=��YY��tʋ5h�S�> t>V�*  �>=Y�Xt"jS�E  �YY��t@VSP�yV  ����uH���> uȋ5h�V�;����%h� �' 3����   Y[_^��5�������%�� �����3�PPPPP�=����U����e� �e� ��VW�N�@��  ��;�t��t	�У��f�E�P�\��E�3E�E���1E��X�1E��E�P�T��M��E�3M�3M�3�;�u�O�@����u��G  ��ȉ��щ�_^��]�U��QW�`���3���tuV��f9t��f9u���f9u�SPPP+�P��FVWPP�8��E���t7P�9  ��Y��t*3�PP�u�SVWPP�8���u	S����Y3�W�d����	W�d�3�[^_��]�U��`�3�t�u��]�]�%��U��d�3��ut��]����]�U��h�3��ut��]����]�U��l�3��u�ut��]����]�U��p�3�t�u�u�u��]��u�u�p�3�@]�U��QV�5����y%���3�3��u�tV�M�Q�Ѓ�zuF�5��3���^����]�VWh������50���h��W��3�h��W�`���3�hȞW�d���3�hԞW�h���3�h��W�l���3�h��W�p���3�h�W�t���3�h �W�x���3�h8�W�|���3�hP�W�����3�hd�W�����3�h��W�����3�h��W�����3�h��W�����3�hȟW�����3����hܟW��3�h��W�����3�h�W�����3�h4�W�����3�hT�W�����3�hh�W�����3�h��W�����3�h��W�����3�h��W�����3�h��W�����3�hȠW�����3�hؠW�����3�h��W�����3�h�W�����3�h�W�����3�h,�W�����3����h<�W��3�h\�W�����3�_���^�U���u�t�]�U���u�x�P�|�]�U��j �l��u�h�]�U��VW3�j �u�u�_  ������u%9��vV�������  Y;5��v������uŋ�_^]�U��SVW�=��3��u�������Y��u#��tV�X����=�����  Y;�v������u�_^��[]���U��VW3��u�u��]  ��YY��u*9Et%9��vV�	������  Y;5��v������uË�_^]�VW�0��0�����t�Ѓ�;�r�_^�VW�8��8�����t�Ѓ�;�r�_^�������������h� d�5    �D$�l$�l$+�SVW��1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q��������U���S�]VW�E� �{�s3=��E�   ����t�O�30�����G�O�30�����E�@f��   �E�E�E�E�C��C�E������   �@�@�L�����E���t{���R  ��M����~   ~h�E�8csm�u(�=L� thL��tZ  ����tj�u�L����U�M��Q  �E�U�9Pth�V����Q  �E�X����tu�f�M��]��Ã���^�����tG�!�E�    ��{�t6h�V�˺�����Q  ����t�O�30��~���W�O�32�~���E�_^[��]ËO�30�~���G�O�30�~���M��֋I�Q  �U���5������t�u��Y��t3�@]�3�]�U��E���]�j��]  Y��tj��]  Y��u�=��uh�   �1   h�   �'   YY�U��M3�;�x�t
@��r�3�]Ë�|�]�U����  ��3ŉE�V�uWV������Y���y  Sj�R]  Y���  j�A]  Y��u�=����   ���   �A  h�h  h ���[  ��3ۅ��1  h  h2�Sf�:������  ��uhL�Vh2��[  ������   h2���[  @Y��<v5h2���[  jh|��E����-2���+�VQ��[  ������   h��h  � �V��Z  ������   Wh  V�Z  ����u}h  h��V�~\  ���Wj��@�����tI���tD3ۋˊO�����f9Ot	A���  r�S������]�P�����P�  YP�����PV���[�M�_3�^�>|����]�SSSSS����������������������7   ���"�.   ��������2��ƅp��������������
�t����
�t�����������������������ݽ`������a���u2����X��������-ʄ���
�t����
�t�������
�t�����������؊�� ����������������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�	]  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�\  ���$��'  �   ��ÍT$�'  R��<$tmf�<$t�I'  =  �?s+��������������=`� ��'  �   ����'  w:�D$��%�� D$u)��   ����-ʄt�����'  ���� u�|$ u����-���   �=`� �J'  �   ����S&  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�9a  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u��`  ���$�&  �   ��ÍT$�=&  R��<$tL�D$f�<$t�-���  �t^�   �uA������=`� �\&  ����   �Y&  �   �u�ԩ�� u�|$ u%   �t����-���   �"�%  ���� uŃ|$ u����-*��   �=`� ��%  ����   ��$  Z�U���uj �u�u�u�   ��]�U��� �e� 3�W�}�jY�9Eu�����    �G�������x�EV�u��t��u������    �#�������S�����M�;�w�E��u�E��E�B   �u�u��u�u�P����������t�M�x�E��  ��E�Pj �
���YY��^_��]�U��} u�i����    謲�����]��uj �5�����]��54����U��E�,��0��4��8�]�j$hP��3����e� �e� 3ۉ]�3��}؋u��Pt��jY+�t"+�t+�t^+�uH�*������}؅�u����b  �E�,��,��^�w\V�Q  YY���E� �V�ƃ�t6��t#Ht�����    �ֱ����E�4��4���E�0��0���E�8��8�3�C�]�P���E܃���   ��uj�D�����tj ��F  Y�e� ��t
��t��u�G`�Eԃg` ��u?�Gd�E��Gd�   ��u-�h��щU̡l��;�}$k��G\�d B�Űh���j � ��M��E������   ��u �wdV�U�Y��u�]��}؅�tj �G  Y�V�U�Y��t
��t��u�EԉG`��u�EЉGd3�������U��U�`�V�u9rtk���E;�r�k�M;�s	9ru���3�^]�U��E��t���8��  uP�+���Y]�U��SVW3���   �;�+���jU�4�P��u�   ����ty�^���~;�~Ѓ�����T�_^[]�U��} t�u����Y��x=�   s	��0�]�3�]�U����3�t3�QQQ�u�u�u�u�u�u��]��u�u�u�u�u�u����YP���]�U��V�u3���t^�MSW�}jA[jZZ+��U�jZZ�f;�rf;�w�� ������f;�rf;Ew�� ����Nt
f��tf;�t�����_+�[^]Ã%H� áD�Vj^��u�   �;�}�ƣD�jP�����@�YY��ujV�5D������@�YY��ujX^�3ҹ����� �R��(�}�@���3�^��_  �=�� t�]  �5@��]����%@� Yø���U��V�u���;�r"���w��+�����P�C  �N �  Y�
�F P���^]�U��E��}��P�qC  �EY�H �  ]ËE�� P���]�U��E���;�r=�w�`���+�����P�D  Y]Ã� P���]�U��M�E��}�`����AP�gD  Y]Ã� P���]�U��E��u�K����    莭�����]Ë@]�U��M���u�&���� 	   �8��x$;��s�������������D��@]������ 	   �4���3�]�jhp������3ۉ]�u���u萻���轻��� 	   �   ����   ;5����   ���������������D8��u
�G����  �jV�^  Y�e� �����D8t�u�uV�^   ������E���� 	   �����  ����}��E������
   ���(�u�}�V�2_  Y��ں�������� 	   �J�������[����U���  �`  ��3ŉE���D��� �E�MV3���8���W3���0�����@���9uu3��  ��u�n���!0蛺���    �ޫ�������  �Ћ���������(���S������$����\$�����t��u+�E�Шu����!0�@����    胫���  ��8����D tjj j P�  ����8��������Y���P  ��(�����$��������D��2  ����3ɋ@l9��   �����P��(�������<�����$��������4�������  9�<���t����  �����0���3�!�8����������4�����,���9M��  ��,���3҉�@���ǅ���
   !�<�������  �3���$�����
���������(���������<���9|8t�D4�E�<����U�j!|8�E�P�Z��P�  Y��tD��0�����,���+�E����  jR��4���P��]  ������  ��,���@��@����&j��,�����4���P��]  �������  ��,���3�@��@���QQj��,����E�Pj��4���PQ������8���<�������  j ��8���Q��$���P�E�P��(��������4������L  ��@�����D����<���9�8����I  9����tK��$�����8���j Pj�E��E�P��(��������4�������   ��8�����  ��D���F��4����   ��t��u3�3�f;������4�������<�����@�������,�����@�����t��uKQ�\  Y��4���f;�uu��9�<���t"jXP��4����h\  Y��4���f;�uOF��D�����@�����,���;U������E  ��(���F���$��������D
4�����D8   �  �����
  ��(���������$����D��u  ��0���3���4������  �]��8�������  3ɍ�������<���+�0���;�sD�
B@�������
��8�����<���u��D����GA������G��8���A��<������  r���$���������+��� ���j PW������P��(��������4���������� ���9� ���|��8�����+�0���;��A�����4�����D�������  ����  j[;���  耵��� 	   �A������  �ʀ���   9u�|  ǅ���
   ����� ��������j+����^;Es3�9����f;����u��D���f�3����f�;�������  rȍ�������<�����$���+�j �� ���PS������P��(��������4�����@�����4����������� �����@���9� ����������<�������0���+�;E�.���������]��8�������  ǅ���
   ����� ��H�����8���+ʋ����;�s;�7������8���f;����uj_f�8����8�����f�0�������  r�3�������VVhU  Q��H���+��+���P��PVh��  �8���@�����4�����<������ ���3ɉ�@���j +��� ���RP���������$���P��(��������4�����t��@���� �����<�����@���;�������@�������<�����4���;��������8�����0���+�@���;�������w���j �� ���R�u��0����4������=����� ���3��G���W�Ʋ��Y�<��0�����(�����$��������D@t	�:u3��趲���    �w����  ����+��[�M�_3�^�$i����]�jh����������u؉u܋}���u�8����  �d���� 	   �   ����   ;=����   �����E�߃��������D��tpW��T  Y�e� �E�����Dt�u�u�uW�g   ������������ 	   謱���  �މu؉]��E������   ���+�}�]܋u�W��U  Y��{����  觱��� 	   �����֋�������U��QQV�uWV�8U  ���Y;�u�u���� 	   �ǋ��D�u�M�Q�u�uP�����u��P�$���Y�Ӌƃ����������d0��E��U�_^��]�U���D�V�   V�M���Y�M�A��t	�I�q��I�A�A�A   �A�a �^]�U��U3�SVAW�����rx��t�������   ��t�����r|��t�������   ��t����j�r[�~�T�t�>��t�����~� t�~���t������Kuҋ��   �   ��A_^[]�U��SV�u3�W���   ��tf=ؾt_�Fx��tX9uT���   ��t9uP�'������   ��U  YY�F|��t9uP�	������   �V  YY�vx�������   ����YY���   ��tD9u@���   -�   P�Ȏ�����   ��   +�P赎�����   +�P觎�����   蜎�������   =X�t9��   uP�V  ���   �s���YYjX���   �E�~��T�t���t�8 uP�H����3�A���YY�E�� t�G���t�8 uP�$���Y�E����H�Eu�V����Y_^[]�U��U����   SV���W�����Jx��t�������   ��t�����J|��t�������   ��t����j�J[�y�T�t�9��t�����y� t�y���t������Kuҋ��   ���   ��1N_^[��]�jh���`����e� �l������x��Npt"�~l t�T����pl��uj �j���Y���n����j�4  Y�e� �5���FlP�!   YY���u��E������   뼋u�j��5  Y�U��W�}��t;�E��t4V�0;�t(W�8�����Y��tV�����> Yu����tV�F���Y��^�3�_]Ã=�� uj��M  Y���   3��U��E-�  t&��t��tHt3�]áP�]áL�]áH�]áD�]�U����M�j �����%`� �E���u�`�   ����,���u�`�   �������u�E��`�   �@�}� t�M��ap���]�U��S�]VWh  3��sWV������{3��{����  �  �{����0�+��7�FIu���  �   �9�AJu�_^[]�U���   ��3ŉE�SV�u������WP�v�İ3ۿ   ����   �È�����@;�r�����������ƅ���� ��Q���;�sƄ���� @;�v�����u�S�v������PW������PjS�Y  S�v������WPW������PW��  S�TX  ��@������S�vWPW������Ph   ��  S�,X  ��$����M�����t�L��������t�L ��������  ���  A;�r��Yj���  ��X+������������� ��w
�L�A �������w��H �A������������  A;�r��M�_^3�[�^a����]�jhИ�����3��u���������x��Opt9wlt�wh��uj �����Y��������j�1  Y�u��wh�u�;5T�t4��t�����u��0�tV�s���Y�T��Gh�5T��u�3�@���E������   둋u�j�"2  Y�jh��8�������E����؉]��<����sh�u�����Y�E;F�h  h   �%���Y�؅��U  ��   �E��ph���3��3S�u�A  YY���}���  �E��Hh�����u�Hh��0�t
Q誈��Y�E��Xh3�@���E��@p��   �x���   j��/  Y�u��C�H��C�L���  �\��ΉM��}f�DKf�MP�A��ΉM��  }�D��(�A��u��   }��  ��0�F��T������u�T�=0�tP����Y�T�3�@���E������   �1�}j�0  Y��#���u��0�tS谇��Y茨���    �3���������U��� ��3ŉE�SV�u�u�6�����Y��uV����Y3��  W3��ϋǉM�9�X���   A��0�M�=�   r����  ��   ����  ��   ��P�������   �E�PS�İ����   h  �FWP������^��3ۉ�  C9]�vO�}� �E�t!�H��t�����LA;�v����8 uߍF��   �@Iu��v�"�������  �^��~3��~����   9=`�tV�����   ����   h  �FWP�]�����kE�0�E���h��E�8 ��t5�A��t+������   s��P�DB�A;�v���9 u΋E�G���E��r�S�^�F   �o�������  �E��Nj��\�_f��Rf��IOu�V�I���Y3�_�M�^3�[�%]����]�U����u�M��V����E�ȋE����   �H% �  �}� t�M��ap���]�U��j �u����YY]������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�3���9d����U���S�]W�}��u��t�E��t�  3���E��t��V�����v�b���j^�0視���X�u�M��#����E�3�9��   ubf�E��   f;�v;��t��tWVS�B���������� *   �����0�}� t�M��ap���^_[��]Å�t��t_��E��t��    �эM�uQVWSj�MQV�p�8��ȅ�t9uu��E��t�������zu���t��tWVS�����艤��j"^�0�͕���o���U��j �u�u�u�u�������]��V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� S��QQ�����U�k�l$���   ��3ŉE��CV�sW���|����Ht+Ht$HtHtHtHHtHuzj��   �nj�
j�j�j_Q�FPW�!  ����uG�K��t��t��t�e����E��F�����]��E��FP�FPQW��|���P�E�P� #  ����|���h��  Q�(  �>YYt�=|� uV蒷��Y��u�6��%  Y�M�_3�^�YY����]��[���U�������$�~$�   ��fD$f%��f��fW�f����fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU��fV�f($������X��\��Y��Y��Y����X��^�f8�f-(��\�fs�?��fs�?�Y�fp�Df50��Y��Y���fW��Y�f\%���Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<����Y��Y��Y��\�fT���X��\��X�f-(��\��X�f8��^�f0�fX������Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(5@�f�f(P�f(%`�fY�f(-����fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT=��f%��f(@��Y�f(P��\�f(`�fp�D�Q�fY�fp�Df��fY�fX�f �fY�����Y�fX�fp�D�Y�fT��fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�P���fD$����fD$�D$���f������fn�fp� f��f��fT�fT��X�fD$�D$���f��f���X�fD$�D$���fW��Xƺ�  �J���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�U������E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z����������������������   s�������������������������   v��������U�������$�~<$�   ���~|$f�f(�fT0�f/X���  �U  f/H�snf/P���  f(�fY�f(�fY�f(- �fY�fX-��fY�fX-��fY�fX-���Y�f(�f���X��Y��\�f�|$�D$�f/@���   f(�fY�f(�fY�f(-��fY�fX-��fY�fX-��fY�fX-��fY�fX-��fY�fX-p�fY�fX-`�fY�fX-P��Y�f(�f���X��Y��\�f�|$�D$��~�fW�f/8�sO�~0��~-��~��X�fs�,f��f~؍@�~,�ȅ�~��\��Y��X(��^�f���   �~��~ ��^�f��~Ÿ��~$���f(�fY�f(�fY�f(- �fY�fX-��fY�fX-��fY�fX-���Y�f(�f���X��Y��\��\��\�fV�f�D$�D$�f/�u�D$�f/`�s�h��h����$�$���D$��h��h��D$��~��~ �fT�f.�z�D$���h���@�ú�  ���T$�ԃ��T$�T$�$��������D$Ð����U�������$�~$�   ��fD$f��f%�f-00f=��B  f���Y�f���-��X�f���\�f(���Y�fɁ�v ����?f(-���p����fY��\��Y���\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-���Y fX5p�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f ��\�fL$�D$��������I ����U�������$�~$�   ��fD$f�f(��f(5`�f(��f(��f��%�  ��@  +�-�<  Ё�   ��(  fY�fX�f(�f\�fY�f(%��fY�f(-��f\�f~��ȃ�?������f\�f(���fY�f(�fY�fX��Y��X�f�fo5@�f��fo5P�f��fs�.fY��X�fV�f��X���~  ��|  w�Y��X�fD$�D$��Ã���|$f�T$f�� f�$�,$����+�fo50�f���  fn�fs�4fV���  fn�fs�4f$�$ft$�D$����f$$�$���$f$�l$��f�����  ���  s'�� t)�Z��   �r��+#��rJw�T$���9��r<��   ��   ��fD$�T$�ԃ��T$���T$�$����fD$����fD$�D$���=  �s1�D$=   �sf ��Y��   �f��Y��   뉋T$=  �w�� u�D$=  �u�������ú�  �V����D$%���=  �@s�fD$�X����fD$�D$��ÍI ƅp����
�u;�����ƅp����2������+  ������a���t������@u��
�t���Ҙ���F  �t2��t��������Ș���^��������- �ƅp����������ݽ`������a���Au����ƅp������-*��
�uS��������
�u�����n�����   ����
�u���u
�t���ƅp����- ���u�
�t��������-������Ș��X��ݽ`������a���u���- �
�t���ƅp�������������- �ƅp����
�u����- �������->��ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���R������ٛ���t�   ø    ���   ��V��t��V���$���$��v��  ���f���t^��t��������������U���������$�\$�   ��fD$f=1f 1fT���fs�,f�� fV�f��%�   ��%�  �Y<���f,����f(4�����  +у�ʁ�   ���  �    �� fn�f��fs����fh1��fs�&f�� fT%1%�   ��%�  �Y���Y,���fX4��fV% 1�X�fT���fs�f�� fh1�\�f=p1%�  ��%�  �Y,���Y��fX4��fT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�fh1f���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%h1fT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f(�(�Y��-��Y�f(�(�X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X 1fY��\ 1fY��\�����f(� )f(5@1fY�fX�fp���Y�fW���?  �X�f���X�f%`1fn��YT$�Y�fs�-fp�Df(=P1�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��XŃ��X��X��X�fD$�D$���fL$f01f~���fT�fs� f~Ɂ�  ���   ��� �  �� �  �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$fT$��  fn�fT01fs�4f��f�1f��fv�f��%�   �� ȁ�   ��r^�� f1f 1�&���f|$fd$f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=1f 1�Y�f~�fs� f~��� tRfT���fT01fs�,f�� fV�%�   ��%�  �Y<���f,����f(4����> �\����Ё������ u��T$��   ��� t1��#��  ��fn�fs� f 1fT$�^ʺ   �  ��#��� ��   ���f1fW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   uefL$fT$��  fn�fT01fs�4f��f��f��fv�f��%�   =�   t#fL$f��% �  �� t��1���1�fL$f��% �  �� �G  ���fL$f��% �  �� �+  ����X��ĺ�  �  fT$f~�fs� f~ҁ����¹    �� �����fx1f�1�Yɺ   �H  fd$fT$f1fW�fT�fv�f��%�   =�   ��   f~��� u fs� f~��  �?��   ��  �u���f1fW�fT�fv�f��%�   =�   uUf��fd$% �  ��  �у� ��   �� tf��%�  =�?  r���f��%�  =�?  s�����1��X��º�  �cf~�fs� f~��������f 1�   �� t:f~�   %���=  �w%r�� w��fD$�D$���f���   ��fD$�T$�ԃ��T$���T$���$�����D$��Ã� ~(=   �<  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X 1���� fY��\ 1fY��\�����f(� )f(5@1fY�fX�fp���Y��X��X�f%`1fnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(=P1�X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� N^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� ������fD$�D$���^�X��Y��Y��X�f��%�  �   =�  ������   �� �������fD$�D$���f�1fn��Y�fs�-fV��   �����   �� tf�1�Y�1�e���f�1�Y��T���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r �ɀ� fn�fs�-��fD$�D$���fd$f�����  ���?  f��3�% �  �� �-����K�����$    ��$    �U��QQ�EQQ�$��4  YY��uJ�EQQ�$�C  �E����YY����Dz+���QQ�U��$�   �E�����YY��DzjX�	3�@���3���]�U���E�  �V3���  ��9Mu:9uu|��������z�����h���   ��������A�E��   ������   9EuB9uu=��������z�������   ������A�Eu�h��   �p�3��F�   ��9Mu-9u��   ���E������A�m����������E{[�����U9Eu]9uuX�EQQ�$�������EYY�ы�����Au�����h���u���������z��u������E��	�M�������^]���U�������$�~$�   ��fD$f��f%�f-00f=��B  f :�Y�f:�-��X�f :�\�f(:�Y�fɁ� v ����?f(-�9��1���fY��\��Y(:�\�fxf����\�fY�f\�f(5�9�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�9�Y fX5�9fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y@:fD$�D$���f0:�Y��\��Y8:fD$�D$����ؔ���U��QQ�E���]��E���]�U��E� tj��t3�@]ètj��tjX]������]�S��QQ�����U�k�l$���   ��3ŉE�V�s �CVP�s�   ����u&�e��P�CP�CP�s�C �sP�E�P�  �s ���s�c����=|� Yu)��t%�CV���\$���\$�C�$�sP�  ��$�P�X  �$��  V��  �CYY�M�3�^��8����]��[�U���S�]V�����t�Etj��  Y����  ��t�Etj��  Y����u  ����   �E��   j�  �EY�   #�tT=   t7=   t;�ub�M������x���{L�H�M�������{,�x��2�M�������z�x���M�������z�h���h���������   ����   �E��   W3���tG�M���������D��   ��EPQQ�$��  �E�� ����E�U���=����}3���G�W��3�����AuB�E���������f�E��E;�})+ȋE��E�t��uG���E��E�t   ��E��m�Iu��E��t���E��3�G��_tj�X  Y�����t�E tj �B  Y���3���^��[��]�U��=|� u%�u�E���T$���\$�$�uj�W  ��$]��$���h��  �u� !   �  �EYY]�U��j �u�u�u�u�u�u�   ��]�U��E3�S3�C�H�EW�  ��H�E�H�M��t�E��  �	X��t�E��  ��H��t�E��  ��H��t�E��  ��H��t�E��  ��H�MV�u�����3A��1A�M����3A��1A�M�����3A��1A�M�����3A��1A��M����3A#�1A�;  ����t�M�I��t�E�H��t�E�H��t�E�H�� t�E	X��   #�t5=   t"=   t;�u)�E��!�M���������M��������E� ���   #�t =   t;�u"�E� ���M�������M�������E�M��3���� 1�E	X �}  t,�E�` �E� �E�X�E	X`�E�]�``�E��XP�:�M�A �����A �E� �E�X�E	X`�M�]�A`�����A`�E��XP�b  �EPjj W�Ȱ�M�At�&��At�&��At�&��At�&��At�&ߋ��������� t/HtHtHu(�   � �%����   ���%����   ��!������� tHtHu!��#�   �	�#�   ��}  ^t�AP���AP�_[]�U��E��t�����w��|��� "   ]���|��� !   ]�U��U�� 3ɋ�9ŀ�t@��|���ń��M��tU�E�E�E�E�E�E��EV�u�E�E h��  �u(�E��E$�u��E��  �E�P��������uV�Y���Y�E�^�h��  �u(��  �u�=����E ����]�U���E������W��Dz	��3��   Vf�u�Ʃ�  u|�M�U���� u��tj�ٿ�������Au3�@�3��EuɉM��y���M�O�Et�f�u�U���  f#�f�u��t� �  f�f�u�Ej QQ�$�1   ���#j Q��Q�$�   ���������  ���  ^�E�8_]�U��QQ�M�E�E�����  %�  ���]��f�M��E���]�U��}  ��Eu��u@]Á}  ��u	��ujX]ËM��  f#�f;�uj���  f;�u�E�� u��tj��3�]�jh������=��|[�E�@tJ�=�� tA�e� �U�.�E� �8  �t�8  �t3��3�@Ëe�%�� �e��U�E������
�࿉E�U�Ͱ���U��Q�}����E���]�U��Q��}��M�E��#Ef#M�f����E�m�E���]�U��QQ�M��t
�-���]���t����-���]�������t
�-���]����t	�������؛�� t���]����]�U��Q��}��E���]�U��V�u��t�U��t	�M��u��y��j^�0��j����^]�W��+���A��tJu�_��u��ty��j"��3���U��V�u�<��� uV�q   Y��uj褠��Y�4������^]�VW�����S���t�tS�H�S�3X���' Y����о|�[�> t�~u�6�H�����о|�_^�jh0�������=�� u����j�i���h�   ����YY�}3�9���u\j����Y����u�x���    3��Bj
����Y�]�9���uSh�  V�5������4����V�xW��Y�E������	   3�@謮���j
�;   Y�VW����h��~uj �>��h�  �6�ߩ��������о|�3�_@^�U��E�4Ű����]����������������SVW�T$�D$�L$URPQQh�Rd�5    ��3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�R'  �   �C�d'  �d�    ��_^[ËL$�A   �   t3�D$�H3���-��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�&  3�3�3�3�3���U��SVWj Rh�SQ�0N  _^[]�U�l$RQ�t$������]� U����u�M��Si���M��yt~�E�Pj�u�m&  ��������   �E�A���}� t�E��`p�����]�U��=(� u�M�P��H��]�j �u����YY]�U����M�SW�u��h���]�   ;�s`�M�yt~�E�PjS��%  �M������   �X����t�}� ���   �t�E��`p�����   �}� t�M��ap����   �E�xt~-�ÍM����EQ��P�����YY��t�Ej�E��]��E� Y��Uu��3�A� *   �]��E� �E�U�j�pjRQ�M�QW���   �E�P��!  ��$��u8E��{����E��`p��o�����u�}� �E�t%�M��ap���U��E���Ѐ}� t�M��ap���_[��]�U��=(� u�M�A���w�� ��]�j �u����YY]���U��W�=����   �}ww�U�����fn��p� ۹   #σ����+�3��of��ft�ft�f��#�uf��#���ǅ�EЃ������Sf��#���3�+�#�I#�[��ǅ�D�_���U��t93���   t�;�Dǅ�t G��   u�fn�f:cG�@�L�B�u�_�ø����#�f��ft �   #Ϻ������f��#�uf��ft@��f����t����뽋}3�������ك��E���8t3�����_��U��UV�uW�z��u�Ps��j^�0�d�����   �} v�M� ��~���3�@9Ew	�s��j"���0S�^�Å�~���t��G�j0Z�@I���U�  ��x�?5|�� 0H�89t�� �>1u�B�S����@PSV�R����3�[_^]�U���,��3ŉE��E�M�SV�uW�u�E�E�E��be���E�3�PWWWWV�E�P�E�P�b.  �؃� �E��t�M��u�E�P��(  YY��u��t��uj���u���tj_�}� t�M܃ap��M���_^3�[�(����]�U���(��3ŉE�SV�u�M�W�u�}��d���E�3�PSSSSV�E�P�E�P��-  �E�E�WP��"  �ȃ�(�E�u��t��uj�
�u��tj[�}� t�M��ap��M���_^3�[�(����]�U��j �u�u�u������]�U��QQ�ESVW�x�   ��P�ϋ �� �  ������ ���  �}���E���t���  t�� <  �%��  �!��u��u�E!P!f�x�X��<  3����M�����������E�]�s���x&�����ʁ���  ����y�}�}��E�s�f�{_^[��]�U���0��3ŉE��ES�]V�E܍EWP�E�P����YY�E�Pj j���uЋ���f���3  �u܉C�E��E��C�E�P�uV������$��u�M���_�s3�^[�&����]�3�PPPPP�va������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��U��M�E������#�V�u�����t$��tj j ��<  YY���n��j^�0�!`�����Q�u��t	��<  ����<  YY3�^]�j����Y������������U��E3�SVW�H<��A�Y�����t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�hP�h� d�    P��SVW��1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�jhp��s���胑���@x��t�e� ���3�@Ëe��E�������\���h�\� �����U��E���]�U���V�u�M���_���E�M���E�L0u3�9Ut�E����   �p#E���t3�B�}� ^t�M��ap���]�U��jj �uj ������]�U��} u�u��K��Y]�V�u��u�u�K��Y3��MS�0��uFV�uj �5���԰�؅�u^9(�t@V�Z���Y��t���v�V�J���Y�.l���    3�[^]��l������P�"l��Y����l������P�
l��Y�����U��V�u��tj�3�X��;Es��k���    3��Q�u��uF3Ƀ��wVj�5�����ȅ�u*�=(� tV謣��Y��uЋE��t�봋E��t�    ��^]�U��VW�}��t�M��t�U��u3�f��Rk��j^�0�\����_^]Ë�f�> t��Iu��t�+��f��Rf��tIu�3���u�f��k��j"�U��V�u��t�U��t�M��u3�f���j��j^�0�+\����^]�W��+��f��If��tJu�3�_��u�f��j��j"��U��Ef���f��u�+E��H]�U��U�MV��u��u9Mu&3��3��t�E��t��u3�f���u��u3�f��Sj��j^�0�[����^]�S��W�����u+��f�3�vf��t%Ou�� +��f��[f��tOtJu��u3�f���_[�{������u�E3�jPf�TA�X�3�f���i��j"�U��E��x!��~��u���������]��i���    ��Z�����]�U���$��3ŉE��ES� �VW�E�3��EV�E��Ӌ��}��Z����E�95���   h   VhB�а����u&����W�j  VVhB�а�����S  h(BW�0����?  P��h4BW���0�P��hDBW���0�P��hXBW���0�P�ӣ���thtBW�0�P�ӣ��}�� ���t�E��tP�ذ9u�tjX�   9u�t�5���j�����;�tO9=�tGP���5��E��ӋM�E��t/��t+�х�t�M�Qj�M�QjP�U��t�E�u�}��    �0��;�t$P�Ӆ�t�Ћ���t��;�tP�Ӆ�tV�Ћ��}�5��Ӆ�tW�u��u�V���3��M�_^3�[�G����]����U�������$�~$�   ��fD$f%0Zf@ZfW�f8Z��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU�QfV�f($��B���X��\��Y��Y��Y����X��^�f=�Yf-�Y�\�fs�?��fs�?�Y�fp�Df5�Y�Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT=�Yfs���f%@Z���\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<��Q�Y�f(�Y�Y��Y��\��X��\��X�f-�Y�\��X�f�Y�^�f�Yf\ՠB���Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5�Yf�f( Zf(%ZfY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=�Yfp�DfT�Y��f%@Z���\��Y��X��Y��\����Y��Y��\��\��X��\�f(�Yfp���\��X�fp���X��Y��X�fp���^�f( Zf(- Zf(ZfY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(�Y�Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�+j��fD$����fD$�D$���f0Zf�Yf�Y�X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$���U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(pZf(�Zf(%�Zf(5�ZfT�fV�fX�f�� %�  f(�P[f(�`_fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f( [f(�f(0[fY�fY�fX�f(@[�Y�f(-�ZfY�f(��ZfT�fX�fX�fY��Y�fX�f(�f�fY˃�f(�f��X��X��X�fD$�D$���fD$f(�Z��� f�� �� wH���t^���  wlfD$f(pZf(�ZfT�fV���� f�� �� t�[ú�  �Of�Z�^�f [�   �4f�Z�Y�������/��������  ���  s:fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$�Lg���D$���fT$fD$f~�fs� f~с��� ��� t���  릍d$ Q�L$+ȃ����Y�J  Q�L$+ȃ����Y�4  jh��訕��3��}�j����Y!}�j^�u�;5D�}S�@�����tD�@�tP�j1  Y���tG�}��|)�@����� P�H��@��4��@>��Y�@��$� F��E������   ���i���Ë}�j�����Y�U��V�u��u	V�   Y�/V�,   Y��t�����F @  tV�h���P�M1  ��YY��3�^]�U��SV�u3ۋF$<uB�F  t9W�>+~��~.W�vV�%���YP薢����;�u�F��y����F��N ���_�N�Ãf �^[]�j�   Y�jh���X���3��}�!}�j����Y!}�3��]�u�;5D���   �@�����t]�@�tWPV����YY�E�   �@����@�t0��uP�����Y���tG�}����u�@tP�����Y���u	E܃e� �   F녋]�}�u�@��4�V����YY��E������   ����t�E��Փ��Ë]�}�j�^���Y�jhؙ�t����}����������4���3�9^u1j
�����Y�]�9^uSh�  �FP�ގ�����F�E������*   ���������������P���3�@�D���Ë}j
�����Y�U��EVW��x`;��sX���������������Dt=�<�t7�=��u3�+�tHtHuQj��Qj��Qj��ܰ������3���_\��� 	   � \���  ���_^]�U��M���u�\���  �2\��� 	   �B��x&;��s�������������Dt�]���[���  ��[��� 	   �6M�����]�U��M���������������P���]�U���SV�u��t�]��t�> u�E��t3�f�3�^[��]�W�u�M��ZN���E����    u�M��t�f�3�G�   �E�P�P�Ŵ��YY��t@�}��t~';_t|%3�9E��P�u�wtVj	�w�4��}���u;_tr.�~ t(�t�13�9E��3�P�u�E�GWVj	�p�4���u��Z������ *   �}� t�M��ap���_�4���U��j �u�u�u�������]�U��Q������u
�..  ������u���  �j �M�Qj�MQP����t�f�E��]����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U��V�u����   �F;�tP�19��Y�F;�tP�9��Y�F;�tP�9��Y�F;�tP��8��Y�F;��tP��8��Y�F ;��tP��8��Y�F$;��tP��8��Y�F8;�tP�8��Y�F<;�tP�8��Y�F@;�tP�8��Y�FD;�tP�}8��Y�FH; �tP�k8��Y�FL;$�tP�Y8��Y^]�U��V�u��tY�;ؾtP�:8��Y�F;ܾtP�(8��Y�F;�tP�8��Y�F0;�tP�8��Y�F4;�tP��7��Y^]�U��V�u���n  �v��7���v��7���v��7���v�7���v�7���v�7���6�7���v �7���v$�7���v(�7���v,�7���v0�7���v4�x7���v�p7���v8�h7���v<�`7����@�v@�U7���vD�M7���vH�E7���vL�=7���vP�57���vT�-7���vX�%7���v\�7���v`�7���vd�7���vh�7���vl��6���vp��6���vt��6���vx��6���v|��6����@���   ��6�����   ��6�����   �6�����   �6�����   �6�����   �6�����   �6�����   �6�����   �w6�����   �l6�����   �a6�����   �V6�����   �K6�����   �@6�����   �56�����   �*6����@���   �6�����   �6�����   �6�����   ��5�����   ��5�����   ��5�����   ��5�����   ��5�����   ��5�����   �5�����   �5�����   �5�����   �5�����   �5����   �5����  �w5����@��  �i5����  �^5����  �S5����  �H5����  �=5����  �25����   �'5����$  �5����(  �5����,  �5����0  ��4����4  ��4����8  ��4����<  ��4����@  ��4����D  ��4����@��H  �4����L  �4����P  �4����T  �4����X  �4����\  �4����`  �t4����^]�U��QQ��3ŉE�SV�uW��~!�E��I�8 t@��u������+�H;ƍp|���M$3���u�E� �@�ȉE$3�9E(j j V�u����   PQ�4��ȉM���u3��q  ~Wj�3�X���rKɍA;�v?�E��E   =   w������܅�t���  �P��3����Y��t	���  ���M���M�3ۅ�t�QSV�uj�u$�4�����   �u�j j VS�u�u賕����������   �E   t,�M ����   ;���   Q�uVS�u�u�y������   ��~Oj�3�X����rC�?�A;�v9�}   =   w�������tg���  �P�3����Y��tR���  ���3���tA�E�WVPS�u�u��������t!3�PP9E uPP��u �uWVP�u$�8���V�B���YS�;���Y�Ǎe�_^[�M�3���	����]�U����u�M��F���u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap���]�U��Q��3ŉE��MSVW3���u�E� �@�ȉEW3�9E W�u���u��   PQ�4��؅�u3��   ~K�����wC��A;�v9�]   =   w��������t����  �P��1����Y��t����  �������t��PWV�w-����SV�u�uj�u�4���t�uPV�u����V�����Y�Ǎe�_^[�M�3������]�U����u�M���D���u �E��u�u�u�u�uP��������}� t�M��ap���]�U��f�M��  f��f#�f;�u-�EQQ�$�t���YYHtHtHt3�@]�j�jX]ø   ]��Ɂ� �  f��u�E�� u�} t��Ƀᐍ��   ]��E��������Dz��Ƀ���A@]���Ɂ������   ]�����U��SVWUj j h(y�u�(  ]_^[��]ËL$�A   �   t2�D$�H�3����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h0yd�5    ��3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y0yu�Q�R9Qu�   �SQ�@��SQ�@��L$�K�C�kUQPXY]Y[� ���U����M�S�u�B���]�C=   w�E苀�   �X�n�ÍM����EQ��P�%���YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�E�PQ�E�P�E�jP�h�������u8E�t�E��`p�3���E�#E�}� t�M��ap�[��]�jh���\������95��t*j����Y�e� Vh���L���YY����E������   �e����j�����Y�U���D��3ŉE��MSVW�A
3ۋ}��% �  �}��E����  �A���?  �E��A�E�����U��E������u%���9\��u@��|��  3��}𫫫j[�  �\��u��}�UܥH�E�j�]ԥ�H����^#�����Uā�  �yI���A+�3�@�uЋ΃����j^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+ȉ]�3�@���EȋD���M�ȉM�;ȋE؋�j�_r;E�s3�A�MԉD��Jx.��t'�D���ˉ]ԍx;��}؋�r��s3�A�MԉD��JyՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA�X���+\�;�}3��}𫫫������;��  +U܍u�UЍ}��¥��������EċEХ%  �yH���@�EЃ���ǉ]��}Ћ�����j �E�X+�j�E�^�T���ϋ���U�#E؋M����T��C�E�;�|ߋEčU���3�j+Ѓ���E�Y;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��E�3��M�@���D����   �����ЅD���9\��uB;�|��v�}̋�j�Y#������  �yO���G�D��+�3�G��ˉ}���}�;��E�j�_r;E�s3�A�D��Jx(��t!�D���ˍx;��}���r��s3�A�D��Jyۃ���MЋUԋ���!D��B;�}�}��΍<�+�3�����`�A���������E؁�  �yI���A�M܋���j �]��׋]�Y+ˉẺM܋T���ˋ���M�#�U��T���M����E��E�@�E�;�|׋u؍U�����j+�3�Y;�|��D����\����Iy������;T���   �`��}�3�������M�   ��������É�  �yI���A����M�j ��X+��]��׉E؋T������#�U��M����MȉT��C�E�;�|ߋu̍U�����j+�3�Y;�|��D����\����Iy�5h�3�5T�C�   �5h��e�����`�������u�����E؁�  �yI���Aj �]������X+ÉM��׉E܋T���ˋ���U�#ǋM����T��F�E���|ߋ}؍U��uȋ���j+�3�Y;�|��D����\����Iy�}�jX+`��ȋE������%   ��d�u���@u
�E�w���� u�7�M���_^3�[� ����]�U���D��3ŉE��MSVW�A
3ۋ}��% �  �}��E����  �A���?  �E��A�E�����U��E������u%���9\��u@��|��  3��}𫫫j[�  �t��u��}�UܥH�E�j�]ԥ�H����^#�����Uā�  �yI���A+�3�@�uЋ΃����j^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+ȉ]�3�@���EȋD���M�ȉM�;ȋE؋�j�_r;E�s3�A�MԉD��Jx.��t'�D���ˉ]ԍx;��}؋�r��s3�A�MԉD��JyՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA�p���+t�;�}3��}𫫫������;��  +U܍u�UЍ}��¥��������EċEХ%  �yH���@�EЃ���ǉ]��}Ћ�����j �E�X+�j�E�^�T���ϋ���U�#E؋M����T��C�E�;�|ߋEčU���3�j+Ѓ���E�Y;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��E�3��M�@���D����   �����ЅD���9\��uB;�|��v�}̋�j�Y#������  �yO���G�D��+�3�G��ˉ}���}�;��E�j�_r;E�s3�A�D��Jx(��t!�D���ˍx;��}���r��s3�A�D��Jyۃ���MЋUԋ���!D��B;�}�}��΍<�+�3�����x�A���������E؁�  �yI���A�M܋���j �]��׋]�Y+ˉẺM܋T���ˋ���M�#�U��T���M����E��E�@�E�;�|׋u؍U�����j+�3�Y;�|��D����\����Iy������;l���   �x��}�3�������M�   ��������É�  �yI���A����M�j ��X+��]��׉E؋T������#�U��M����MȉT��C�E�;�|ߋu̍U�����j+�3�Y;�|��D����\����Iy�5��3�5l�C�   �5���e�����x�������u�����E؁�  �yI���Aj �]������X+ÉM��׉E܋T���ˋ���U�#ǋM����T��F�E���|ߋ}؍U��uȋ���j+�3�Y;�|��D����\����Iy�}�jX+x��ȋE������%   ��|�u���@u
�E�w���� u�7�M���_^3�[������]�U���   ��3ŉE��E�E��E�E�3�S3�@V�E���É]�W�}��]��]��]��]��]�9E$u��C���    �5��3��  �U�ʉM��
�� t��	t
��
t��uB��
B�M����{  �$����A�<wjXJ�݋E$� ���   � :ujX������+tHHt����  3�@�j� �  X�M��jX�]��3�@�E��A�<v��E$� ���   � :uj묀�+t+��-t&��0t���C�:  ��E~��d���)  j�|���Jj�t����A�<�P����E$� ���   � :�R�����0�c����U���  3�@�E���0|*�E��u���9��s	��0@�G�F�
B��0}�u���E��E$� ���   � :�I�����+�t�����-�k����E���3�@�E��E��E���u��0u�E��
HB��0t��E��E���0|%�u���9��s��0@�GN�
B��0}�u���E���+������-������C~��E�������d�������J�	  3���0@�E���	����j�/����B��E��A�<wj	��������+t"HHt�������j����j���X�M������j����3�@�E���
B��0t���1����   몍A�<v���0�9] t"�B��E�����+t�HH�q����M��jX�z���j
XJ��
�m����H3���@�E����93k�
�u������P  �
B�M���0}���M��Q  ���9�
B��0}�J�E��M���M�����  ��v�E�<|���E��M�OjAX�M���M�����  O8u
HAO8t��M��M�QP�E�P�
  �M�����y��u��E���uu�E���u+u��P  �J  �������/  �����`���  y
����ރ�`9]��  3�f�E���  �ƃ�T���U��u�����  k�� �  ʉM�f9r��}��M��M�����M��y
�U΋�3]�% �  �]ԉE���  #Љ]�#��]܍���  �u�f;��I  f;��@  ���  f;��2  ��?  f;�w�]��7  f��u$F�E�����u�u�}� u�}� u3�f�E��  f��uF�A����u�u	9Yu9t�j�ÍU�_�E��}��}���~X�uč4F�A�E���E��E��M��]�� �ȉM�J�;J�r;M�s3�@��E��J���tf��m���O����M��}��E���@O�E��}�����u��U܁��  �}ԉU�f��~;��x2�E؋�����������U��E�Ҹ��  �}����U��U�f���f��i���  �f��y]�]��������E���E�tC�M؋����M��m�	E��E���������M��U܉E؉}�u�j �ۉU�[tf��3�Gf�f�Eԋ}��f�EԺ �  f;�w���� �� � u@�Eփ��u4�Eډ]փ��u f�E޹��  �]�f;�uf�U�F�f@f�E��@�EڋM��@�E֋M��U���  f;�r3��]�f9E��]���H%   � ���E��:f�E�u�f�EċE؉EƉM�f�u�� 3�f9E���H%   � ���Ẻ]ȉ]ċU��u��������E��MċUƋu����23��ˋË�Ӎ_�#��  �   �j��ˋË����Ë�j�ˋ�[�}�E�f�G
��f��W�w�M�_^3�[�.�����]�Ć�p����������C�8��U���   ��3ŉE��U3�S�]��  V� �  �]�#��E������uA#��E������E����?�U��E�Wf��t�C-��C �}f��u:����   9}��   3��Kf�� �  f;�����$ �C��f�C0 ��  f;���   �E�   �f��M;�u��t�   @uh�k�Gf�}� t=   �u��u0h l�;�u%��u!hl�CjP����������  �C�hl�CjP����������  �C3��G  �֋�������3ۉ}濈���`f�u��E�   �H�E���  k�Mi�M  �E��?  ������ȋE�E�3�f�E����؉M��E����/  y�ؿ����`�E����  �u��U�u��}���T�}�����  k�� �  ωM�f9r��}čMĉM�����M��y
� �  �E�}����  1E�%�  !u��E�ǉ}�N���E�f;Ƌu��]��]��]�]��}��X  ��  f9M��M��F  f;}��<  f;}�w�]��E  f��u G�E�����}�u��u��u3�f�E��-  f�}� uG�A����}�u	9Yu9t�j�ÍU�^��|����u��u���~r�u��F�q��x����u��u��M��8����B��]��8;ȉM���r;�s3�A��M��B���tf���x����M�������x���N�M�����M��u���|�����@N��|����u����q����}��E����  �u��E�f��~;��x2�E�֋���������E�E���u�����  ��E��E�f���f��q���  �f��ye�]�����3�����E��}�B�}��U�tG�M�����M��m�	E��E���������M��]��E�u�u�j �]����}�[tf��f�f�E��u��f�E� �  f;�w���� �� � u@�E���u4�E��]���u f�E����  �]�f;�uf�M�G�f@f�E��@�E��M��@�E�M���  f;�s f�E�}�f�E��E�E�u��M�U�f�}��!3�f9E���H%   � ���E��Ӊu��U�u��}��E���������M���U�u��E��?  ��f;���  A�]��M��ȋEڋ�3��]��� �  �]�}���  #ǉ]�#ωE������  �}�f;��@  �E�f;E��3  f;}��)  f;}�w�]��2  f��u G�E�����}�u��u��u3�f�E��  f��uG�E�����}�u�}� u�}� t��ӍM�j�U�X����~X�}��E؍<W�E��}����ЋA��]��<;�r;�s3�@��E��y���tf��}��E������}�N�E�����U��E���BH�U��E�����}��u����  f����   �]��]���x,�E�Ӌ���������E�۸��  �]����u�f��Љ]��U�j [f��~[f�M� �  f;�w���� �� � ��   �E�����   �E��]�����   f�E����  �]�f;�u|� �  Gf�E��|�U���  �f��y���������E��}��}��E�tG�]�Ƌ��������������M��]�U�u�j ���u��}�[�M���3�f��@f�f�M��U��<���f@f�E��@�E��u��@�E��  f;�s f�E�}�f�E��E�E�u�U�u�f�}��3�f9E���H%   � ���E����E�M��E��}f�t6���}���/3�f�� �  f9E�����$ �A3�@�A�A0�Y�  �}�jX;�~�E��}������?  3�j�}�f�E�]�_�ʋ���������Љu��]�Ou�}��]��U�u�j [��y7�߁��   ~-�]����������������O�]�u����]�3ۉU�u��u��E�@�E��~�}��ωM�����   �u��ʍ}����ҥ��}������ЋE��4 ��������������E��8�M�;�r;�s�B��;�r��s3�A�ɋЋM�tF�Eȍ<;�r;�sFű��U�������U��U��?����6�U���M��E���0�]�A�E�H�M��E���~�E�E��>����u��}��A���<5|E�	�99u�0I;�s�;�sAf���E�*Ȁ��H�Ɉ\3�@�M�_^3�[�p�����]À90uI;�s�;�s̋M�3�f�� �  f9E�����$ �A3�@�A�0����3�SSSSS��#���U��M3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tƋѻ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t;�u �  ]Ã�@]�@�  ]�U�����}�f�E�3ɨtjY�t���t���t��� t���t��   SV��   ��W�   #�t&��   t��   t;�u��   �
����   ��   t;�u��   ���   ���   ��t��   �}���E��#�#��;���   V�?  ��Y�E��m���}��E�3��tj^�t���t���t��� t���t��   �Ћ�#�t*��   t��   t;�u��   ���   ���   ��   t��   u��   ���   �   ��t��   �=����  ���]�E�3Ʉ�yjY�   t���   t���   t����t���   t��   �л `  #�t*��    t�� @  t;�u��   ���   ���   j@%@�  [+�t-�  t+�u��   ���   ���   ��#}��#��;���   P�$���P�E�Դ��YY�]�E3Ʉ�yjY�   t���   t���   t���   t���   t��   �п `  #�t*��    t�� @  t;�u��   ���   ���   %@�  +�t-�  t+�u��   ���   ���   ���3Ʃ t��   ������_^[��]�U��M3���t@��t����t����t����t�� ��   t��V�Ѿ   W�   #�t#��   t;�t;�u   �   �   �с�   t��   u���_^��   t   ]�U��V�uW�����u�>.���    �����E�F�t9V�t���V���   V�q��P�  ����y�����~ t�v����f Y�f ��_^]�jh���c������}�3��u������u��-���    ������d����F@t�f ��V�lp��Y�e� V�?���Y���}��E������   �ǋu�}�V�p��Y�jh8��c��3��u�}���u�Q-��� 	   �   ����   ;=����   �����E��߃��������D��trW����Y�u��E������Dt(W����YP����u�����u��t�,���0��,��� 	   ����u��E������
   ���!�}�u�W����Y��,��� 	   ���������b��á�����t���tP���3�PPjPjh   @hl������U���S�]3ҸN@  VW�E���S�S9U�<  �ʉU�M�U��U�}�����ҥ���u�΋}��������������������E����s{3ɉE;�r;E�s3�A���t��3ɍp;�r��s3�A�s��tG�{�U�3���M�;�r;�s3�@�K��tG�{�U�u��}���e� �������E���s�{� �u�}��E��M�;�r;�s3�@��E����t$��3ҍp�u;�r��s3�B�s��tG�}��{�EH�s�E�{�E��������N@  3�9Su.�S������������E�����  ��E���tۉS�s�S�� �  u4�;�s�ǋ��������E�����  ��E��� �  tى;�s�S_^f�C
[��]�jhX��`��3ۉ]�u���u�*����K*��� 	   �   ����   ;5��s{���������������D8��u
��)���  �ZV����Y�e� �����D8tV�T   Y�����)��� 	   ����}��E������
   ���(�u�}�V�����Y��|)����)��� 	   ���������_���U��VW�}W�=���Y���tP�����u	���   u��u�@Dtj����j���	���YY;�tW�����YP����u
�����3�W�Y���Y�σ����������D9 ��tV��(��Y����3�_^]�U��V�u�F�t �Ft�v�����f����3�Y��F�F^]�������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �������������%��%̰���̃=�� uK�����t�D�Q�@<�@�Ѓ����    V�5����t���0���V�*��������    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           � �� � � 4� D� P� \� x� �� �� �� �� Ҝ � �� �  � .� F� X� n� �� �� �� ҝ � � &� N� V� j� ~� �� �� �� �� Ğ О � � � � 2� B� T� h� z� �� �� �� �� �� ̟ ڟ �  � � "� 6� D�                   ���*�n�        �z���                    ��DT       O   xl xT     ��DT          �l �T    ��������       ����   ���������������N                     ���������������������������C-DT�!	@-DT�!�?       ����       ����       ����                     ������������       ����       ����       ����         ����    �����������������m�� ���� �� �0�@�`�    0   .   -   ||----------------------------------------  ||  (c) 2012-2014 - Christopher Montesano   ||  http://www.cmstuff.com   v  ||      ||    build date:   �n� 0���P^`�p�� ��� �� ����GP�gui_icons.tif   gui res lo�� �� �`�`� ������ ���6�6�� �6�6�6`��[���7�7�7 �   %  �o�� �]`� �I������e:\repos\cmnodes\src\source\customgui\cmcustomguireal.h CM_REAL_GUI cmRealGUI   p��  �0�@�P�`�p����������������� ���� ��e:\repos\cmnodes\src\source\prefsdialog\cm_prefs.h  Prefs_cm    cmStuff �p�� `�0�@�P�`�p�����������p���`� ������e:\repos\cmnodes\src\source\prefsdialog\cmnodes_prefs.h �pP� P~`~@�P�`�p����������������� ��e:\repos\cmnodes\src\source\nodes\cmnodetree.h  Dq� ���I`������ ����J���������� ��@P`p�������cmNodeTreeRoot  cmNodeBaseRoot  0123456789  StartUndo 11    AddUndo 13  EndUndo 11  AddUndo 14  AddUndo 15  AddUndo 16  AddUndo 17  AddUndo 18  AddUndo 19  e:\repos\cmnodes\src\source\scenehook\cmnodeforest.h    �q �  [�\@�P�`]_�������������\�\ ��`��-���`�� {�g�c�b�fe:\repos\cmnodes\src\source\nodes\node_types\cmnodeoutput.h input   (r0� ���\@�P�0�_�������������\�\ ��`�����`���y0e�cpbx ^ ;AddUndo 20  AddUndo 21  StartUndo 14    EndUndo 14  color   diffusion   luminance   transparency    reflection  environment bump    normal  alpha   specular    displacement    |r�� `��\@�P�`]_�������������\�\ ��0��B��_�b�| e�b���fe:\repos\cmnodes\src\source\nodes\node_types\cmnodeinput.h  �rО `��\@�P�`]_�������������\�\ ��0�p���_�b�| e�b���f$s� p��\@�P�`]_�������������\�\ ����p;��p^�bP{�g�b�b�fe:\repos\cmnodes\src\source\nodes\node_types\cmnodechannels.h   xs�� К�\@�P�`]_������������W�\ ��������p^�b w�d�b`b�finputA  inputB  �s@�  ��\@�P�`]_�������������\p� ��P�@���p^�by�f�b�b�fNormal  Darken  Multiply    Color Burn  Linear Burn Darker Color    Lighten Screen  Color Dodge Linear Dodge    Lighter Color   Overlay Soft Light  Hard Light  Vivid Light Linear Light    Pin Light   Hard Mix    Difference  Exclusion   Subtract    Divide  Hue Saturation  Color   Luminosity  Levr    Grain Extract   Grain Merge mask     t`�  ��\@�P�`]_�������������\�� ��p�����_�by�f�b�b�fe:\repos\cmnodes\src\source\nodes\node_types\cmnodeadjust.h Add Minimum Maximum tt�� ���\@�P�`]_�������������V�\ �� ������_�b�x�d0c`b�f�tП ���\@�P�`]_�������������\�\ ��p� ����_�b�x�d0c`b�fup� @��\@�P�`]_�������������\�\ ����p���_�b�x�d0c`b�fpu@�  ��\@�P�`]_�������������\�� ��P������_�bP{�g�b�b�fLinear -> Linear    Linear  HSV HSL sRGB     ->     �u�� @��\@�P�`]_������������ X�\ �����	���_�b�x�d0c`b�fv � ���\@�P�`]_�������������\�\ ������P��_�b {�g�b�b�flv � ���\@�P�`]_�������������\�\ ��`�����_�b�x�d0c`b�f�v � ���\@�P�`]_�������������\�\ ���� F��P`�bP{�g�b�b�fe:\repos\cmnodes\src\source\nodes\node_types\cmnodeeffects.h    w�� 0��\@�P�`]_�������������\�\ �� �����P`�bx�f�b�b�fsource  displace    hw�� ���\@�P�`]_�������������\�\ ����p��P`�b�x�d0c`b�f�w�� Ч�\@�P�`]_�������������\�\ �����$��P`�b�x�d0c`b�fxp� ���\@�P�`]_�������������U�\ ��б���P`�b�x�d0c`b�fdx�� 0��\@�P�`]_�������������\�\ ��@�P��P`�b {�g0c�b�f�x0� ��\@�P�`]_�������������W�\ ��@�����P`�b�x�d0c`b�fy�� ��\@�P�`]_�������������X�\ �������P`�b {�g�b�b�f`yТ ���\@�P�`�_������������ Y�� ��������a�by e�b���fFacing Ratio    UV Coordinates  Camera Distance Normals (Object)    Normals (World) Normals (Camera)    Object Color    Normal Direction    e:\repos\cmnodes\src\source\nodes\node_types\cmnodeutility.h    �y@� ��\@�P�`]_�������������\�\ ��`��<���a�b�w�g�b�b�fz`� Н�\@�P�`]_�������������\�\ �� ������a�b�w e�b���f\zp� ���\@�P�`]_�������������\�� ����`B���a�b�{�g�c�b�finput 0 input   �z�� ���\@�P�`�_������������ [�\ �����3���a�b�| e�b���f{��  [�\@�P�`]_�������������\�\ ��`��(���a�bP{�gpc�b�fX{ � `��\@�P�`]_�������������\�\ ��������a�bpw�g�b�b�f�{@� ��\@�P�`]_�������������\�\ ��0�����a�b�| e�b���f |�  [�\@�P�`]_�������������\�\ ��`�`C���a�b�| h d�b�ftile    T|� ��\@�P�`]_�������������\�\ ���� 9���a�b�| e�b���f�|� ���\@�P�`]_�������������\�\ ����`)���a�b {�g�b�b�f�|p� ���\@�P�`]_�������������\�\ ����P����a�b v@d�bpb�fcontrol P}P�  ��\@�P�`]_�������������Z�\ ����p.���a�b {�g�b�b�f�}��  ��\@�P�0�_���������M���\�\ ��`����0b�� ~Ph�c�bx ^ <AddUndo 22  AddUndo 23  StartUndo 15    EndUndo 15  e:\repos\cmnodes\src\source\nodes\node_types\cmnodevray.h   matte opacity   matte alpha material weight luminosity color    luminosity dirt luminosity occulded luminosity unocculded   luminosity transparency flakes color    flakes glossiness   flakes orientation  reflection color    reflection transparency specular1 color specular1 transparency  specular1 hilight glossiness    specular1 reflection glossiness specular1 anisotropy    specular1 anisotropy rotation   specular1 reflectance 90 degree specular1 reflectance 0 degree  specular2 color specular2 transparency  specular2 hilight glossiness    specular2 reflection glossiness specular2 anisotropy    specular2 anisotropy rotation   specular2 reflectance 90 degree specular2 reflectance 0 degree  specular3 color specular3 transparency  specular3 hilight glossiness    specular3 reflection glossiness specular3 anisotropy    specular3 anisotropy rotation   specular3 reflectance 90 degree specular3 reflectance 0 degree  specular4 color specular4 transparency  specular4 hilight glossiness    specular4 reflection glossiness specular4 anisotropy    specular4 anisotropy rotation   specular4 reflectance 90 degree specular4 reflectance 0 degree  specular5 color specular5 transparency  specular5 hilight glossiness    specular5 reflection glossiness specular5 anisotropy    specular5 anisotropy rotation   specular5 reflectance 90 degree specular5 reflectance 0 degree  diffuse1 color  diffuse1 dirt   diffuse1 occulded   diffuse1 unocculded diffuse1 transparency   diffuse1 roughness  diffuse2 color  diffuse2 dirt   diffuse2 occulded   diffuse2 unocculded diffuse2 transparency   diffuse2 roughness  refraction color    refraction glossiness   refraction translucency sss overall color   sss color   sss scatter color   sss scatter radius  AddUndo 2   �}�� �=�� ��� �0�@�`�e:\repos\cmnodes\src\source\command\cmnode_commands.h   cut.tif #$  H~�� `=�� ��� �0�@�`�copy.tif    �~�� @>�� ��� �0�@�`�paste.tif   �~�� �=�� ��� �0�@�`�delete.tif  8�� �>�� ��� �0�@�`�select_all.tif  ��� �=�� ��� �0�@�`�deselect_all.tif    ��� �=�� ��� �0�@�`�disconnect.tif  (���  >�� ��� �0�@�`�frame_selected.tif  x��� `>�� ��� �0�@�`�preferences.tif Ȁ��  =�� ��� �0�@�`�add_tree.tif    ��� �>�� ��� �0�@�`�tree_menu.tif   h���  >�� ��� �0�@�`�node_menu.tif   ����  ?�� ��� �0�@�`�zoom_in.tif ���  ?�� ��� �0�@�`�zoom_out.tif    X��� �>�� ��� �0�@�`�zoom_100.tif    ���� �>�� ��� �0�@�`�reset_view.tif  ���� @=�� ��� �0�@�`�calc_preview.tif    03  04  05  06  #$07--  08  09  10  11  #$12--  13  #$14--  15  16  17  #$18--  19  20  21  22  23  H���  C�� ��� �0�@�`� node   Create  node_solid_color.tif    ���� �C�� ��� �0�@�`�node_texture.tif    ��� �?�� ��� �0�@�`�node_clamp.tif  8��� �?�� ��� �0�@�`�node_colorspace.tif ����  @�� ��� �0�@�`�node_curves.tif ؄��  A�� ��� �0�@�`�node_filter.tif (��� @A�� ��� �0�@�`�node_grade.tif  x���  B�� ��� �0�@�`�node_math.tif   ȅ�� @?�� ��� �0�@�`�node_blend.tif  ���  @�� ��� �0�@�`�node_copy.tif   h���  C�� ��� �0�@�`�node_shuffle.tif    ���� `?�� ��� �0�@�`�node_blur.tif   ��� `@�� ��� �0�@�`�node_dirblur.tif    X��� �@�� ��� �0�@�`�node_distort.tif    ���� �@�� ��� �0�@�`�node_edge_detect.tif    ���� �@�� ��� �0�@�`�node_emboss.tif H���  B�� ��� �0�@�`�node_matrix.tif ���� `B�� ��� �0�@�`�node_normal_map.tif ��� �C�� ��� �0�@�`�node_transform.tif  8��� �B�� ��� �0�@�`�node_output.tif ���� �A�� ��� �0�@�`�node_material.tif   ؉�� �?�� ��� �0�@�`�node_colorize.tif   (��� �A�� ��� �0�@�`�node_info.tif   x��� `A�� ��� �0�@�`�node_highpass.tif   Ȋ�� `C�� ��� �0�@�`�node_switch.tif ��� �A�� ��� �0�@�`�node_invert.tif h��� @C�� ��� �0�@�`�node_specular.tif   ���� �C�� ��� �0�@�`�node_vrayadvanced.tif   ��� �@�� ��� �0�@�`�node_distance.tif   X��� �B�� ��� �0�@�`�node_reflection.tif ���� @B�� ��� �0�@�`�node_noop.tif   ���� @@�� ��� �0�@�`�node_diffuse.tif    H���  A�� ��� �0�@�`�node_fresnel.tif    ���� �C�� ��� �0�@�`�node_tiler.tif  ��� �B�� ��� �0�@�`�node_shadow.tif 8��� �?�� ��� �0�@�`�node_condition.tif  ���� �B�� ��� �0�@�`�node_projector.tif  ؎�� �A�� ��� �0�@�`�node_input.tif  ?   Are you sure you want to delete bookmark     has been saved.    Bookmark    d��� 0D�� � � �0�@�`�Tree Bookmark 01    e:\repos\cmnodes\src\source\command\cmtree_bookmark_commands.h  tree_bookmark.tif   ���� 0D�� � � �0�@�`�Tree Bookmark 02    ��� 0D�� � � �0�@�`�Tree Bookmark 03    `��� 0D�� � � �0�@�`�Tree Bookmark 04    ���� 0D�� � � �0�@�`�Tree Bookmark 05    ��� 0D�� � � �0�@�`�Tree Bookmark 06    \��� 0D�� � � �0�@�`�Tree Bookmark 07    ���� 0D�� � � �0�@�`�Tree Bookmark 08    ��� 0D�� � � �0�@�`�Tree Bookmark 09    X��� 0D�� � � �0�@�`�Tree Bookmark 10    0,0 %.0f,%.0f   %.2f    ��P� 0���P���p������ С �Cut Copy    Paste   Delete  Disconnect  Calculate Previews  StartUndo 10    AddUndo 3   AddUndo 4   EndUndo 10  New Tree    StartUndo 2 AddUndo 5   AddUndo 6   EndUndo 2   Error: Could not initialize copy operation  AddUndo 7   cmNodeMat   cmNodeVrayAdv   StartUndo 3 AddUndo 8   EndUndo 3   Error: Could not initialize paste operation StartUndo 4 AddUndo 10  AddUndo 11  AddUndo 12  AddUndo 28  EndUndo 4   unknown StartUndo 5 EndUndo 5   StartUndo 6 EndUndo 6   StartUndo 7 EndUndo 7   StartUndo 8 EndUndo 8   No tree selected    StartUndo 9 EndUndo 9   Add Tree... &c& �� �  � �b�� p���������� Edit    View    Nodes   Bookmark    cmNodeEditor    D��  D�� ��� �y@�`��� � �� � �  � ��У����File    New...  Load... Save... Save All... Copy All    Delete...   Rename...   load    selection   StartUndo 13    AddUndo 25  AddUndo 26  AddUndo 27  EndUndo 13  Are you sure you want to delete     cmtree  Load    Save    cmTreeManager   ��� @G�� ��� �0y@�`�0�`� �� ���cmUpdateNodeThread  e:\repos\cmnodes\src\source\utility\cmbghandler.h   ���� �v 0�@�P��v  z ������������@y �� �� Pw �x �x p����e:\repos\cmnodes\src\source\shader\cmnodeshader.h   Could not find string resource for node     Could not find string resource for category      description    Failed to register  nbase.tif   Node limit exceeded Scmnodeforest   Failed to register cmNodeForest description cmNodes Failed to register cmNodeForest cmNodeTree  Failed to register cmNodeTree   Nbase   Ncolor  Ntexture    Nclamp  Ncolorize   Ncolorspace Ncurves Nfilter Ngrade  Ninvert Nmath   Nblend  Ncopy   Nshuffle    Nblur   Ndirblur    Ndistort    Nedgedetect Nemboss Nhighpass   Nmatrix Ntransform  Noutput Nmaterial   Nvrayadvanced   Ncondition  Ndiffuse    Ndistance   Nfresnel    Ninfo   Nnoop   Nnormalmap  Nprojector  Nreflection Nshadow Nspecular   Nswitch Ntiler  e:\repos\cmnodes\src\source\utility\cmnoderegister.h    #$00cmNodeEditor    Failed to register cmNodeEditor #$01cmTreeManager   Failed to register cmTreeManager    #$02--  cmNode  Failed to register AM Hook  xcmnodeshader   cmNodeShader    prefs_cmnodes   e:\repos\cmnodes\src\source\main.cpp     R14    1001;   1002;   1003;   1004;   1005;   1006;   1007;   Component Failure:  Shaders Cinema4D            ���ư>-C��6?{�G�zt?#���?�������?)\���(�?]m���{�?�������?�v��/�?333333�?
ףp=
�?�������?���z6�?      �?�Q����?���(\��?�A`��"�?333333�?UUUUUU�?�������?]t�E�?      �?�p=
ף�?�(\����?bX9���?333333�?�,C���?      �?�������?ffffff�?      �?�z�G��?�������?       @333333@      @      @-DT�!	@      @      @-DT�!@       @      "@ףp=
�)@      4@      >@      Y@     �b@     �f@     �o@     @@     @�@������      �      �333333�      �?              �?{�G�zt?�������?�������?�������?�������?333333�?333333�?�(\����?��(\���?�������?�������?      �?      �?��Q���?      �?333333�?333333�?      �?      �?333333�?333333�?���Q��?)\���(�?
ףp=
�?�������?)\���(�?���Q��?      �?      �?�������?�������?ףp=
��?333333�?�G�z��?)\���(�?              �?{�G�zt?      �?�������?      �?      �?      �?      Y@      Y@��������������������������       �       ����������������������N���������������C-DT�!	@-DT�!�?��v [�\@�P�`]_�������������\�\ ���a�c0d�d0e@e�e�e�f�foutput  CopyTo - Update StartUndo 1 AddUndo 1   EndUndo 1   TRUE    FALSE   SetNodeDirty:            �V@      �?�������?�������?      �?      �?�������?�������?      �?�������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?�p��������N���������������C-DT�!	@-DT�!�?c:\program files\maxon\cinema 4d r14\resource\_api\c4d_file.cpp �������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?c:\program files\maxon\cinema 4d r14\resource\_api\c4d_basebitmap.cpp   c:\program files\maxon\cinema 4d r14\resource\_api\c4d_misc\datastructures\basearray.h  ,�����*�*�    �������N���������������C-DT�!	@-DT�!�?h�N0�@�P�`�p������� ��T�`N@�P�`�p���������|�`N@�P�`�p�������@0@�`N@�P�`�p�������5ȕ`N@�P�`�p�������@6�6�6�6�6�6�6 77�7�7�7�7c:\program files\maxon\cinema 4d r14\resource\_api\c4d_gui.cpp  ~   Progress Thread 0%  %       ��������������N���������������C-DT�!	@-DT�!�?�h㈵��>����MbP?
ףp=
�?-DT�!�?      @      N@      ^@      n@     �v@      �A-DT�!��       �                -DT�!�?              �A        -DT�!���������N���������������C-DT�!	@-DT�!�?c:\program files\maxon\cinema 4d r14\resource\_api\c4d_general.h       %s      �������N���������������C-DT�!	@-DT�!�?ܕ@� �    c:\program files\maxon\cinema 4d r14\resource\_api\c4d_baseobject.cpp   �������N���������������C-DT�!	@-DT�!�?$��0�l�� c:\program files\maxon\cinema 4d r14\resource\_api\c4d_resource.cpp #   M_EDITOR        �������N���������������C-DT�!	@-DT�!�?����  �0�@�P�`�p����������������� ���� ���������N���������������C-DT�!	@-DT�!�?c:\program files\maxon\cinema 4d r14\resource\_api\c4d_pmain.cpp        c:\program files\maxon\cinema 4d r14\resource\_api\c4d_basetime.cpp        ����A  4&�kC �Ngm��C  4&�k�c:\program files\maxon\cinema 4d r14\resource\_api\c4d_libs\lib_ngon.cpp        fmod         �������T�����������������������      8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7      �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC                                            �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               �       �      ��      ������    ����    ��      ��            8C      8C      0<      0<��+eGW@��+eGW@  ��B.�?  ��B.�?:;����=:;����=�ѱt�?Z�fUUU�?���&WU�?{������?                Mu�{�<`�w>�,  �g5RҌ<t�ӰY  a��aN�`<țuE�  l{�]���<��lX�  ќ/p=�><���2��  ؼcnQ�<P[� {8�&TŤ<�-���B �?RbSQ�<zQ}<�r �S?���<u�o�[� _/:>��<��h1�� �æDAo�<֌b�; �������<8bunz8 ���+G�<�|�eEk 1�	m���<����� �
r�7�<䦅� ���MuM�<�1
� J��]9ݏ<�d�< )}̌/�<ʩ:7�q �^�s)ҧ<���4ۧ mL*�H��<"4L�� ��%F��<).�!
 ��`�cC<-�a`N y����n<�<���� ��z�ΐv<'*6�ڿ 	*(�̃�<�,�v�� ���	�<�O�V+4 ���5�<�'�6Go 	T��c�<)TH�� 5�d+�2�<H!�o� 
���<�U:�~$ �s ��<$"U�8b qU�M��<�;f�� �GΆ�+�<.e<�� �o � �<s_��u ���"a�<�gBV�_ ��F�D�<��s� Ul֫��e<bN�6�� �g�����<�L��% ���<�D��h ����/��<۠*B� D_�Y��{<6w��� <(��`�<��Ͱ77	 �b� ��<ONޟ�}	 'Α+��q<�𣂑�	 �.�X4m�<d�]{f
 ����|'�<\%>�U
 �Zsn�i�<��yUk�
 �3˒w�<��Z���
 �-�f$�<�O��3 ���.�<F^��v ��_
��t<��K�� ��0�ns<�R�ݛ �Y	я��<K�W.�g h�l,kg<i��� � ���6	p�<{�J- �=���t<����X ����PZ�<�2�� ��Js��<^�{3�� ӈ:`�t<�?��.P &I	�'o�<ِ����  �A�Î<'Za�� ��1�d�<@En[vP �͑M;�w<ؐ����       �?       �9��B.�@  ׽2b      �        �������         0<  0<�dW�dW      �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �      �?      �?3      3                      �                     �              �?      �?3      3            �      0C       �       ��              ̖���          8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �        ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=(null)  ( n u l l )            EEE50 P    ( 8PX 700WP        `h````  xpxxxx          x���    �������             ��      �@      �               ���5�h!����?      �?            �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��log log10   exp pow asin    acos    exp10   atan    ceil    floor   modf    sin cos tan sqrt       �U��?�wB%�K�=      �?   �[��?(�6N�g�=      �?   $�?V�`t� >      �?   ��տ?��2n{a>      �?   ����?��M��=      �?   H{��?{4�r>      �?   Pא�?"�"�>      �?   �u[�?��*��>      �?   ����?G�0��_(>      �?   4wb�?��i^^?(>      �?   ��0�?p3���>      �?   @��?F��M>      �?   8M��?�B�V��>      �?   ��d�?}B��a.>      �?   ȴ�?d�����>      �?   g��?�ߊ��>      �?   �@�?�f\���*>      �?   �~e�?�-��f>      �?   �]%�?D	�G��?>      �?   ���?�\����>>      �?   X���?�1��#>      �?   �E�?��h��>      �?   �?��?�ⳇ��>      �?   ����?�$	�49>      �?   x�8�?k���0H<>      �?   ����?r��ش8>      �?   8fm�?�"m>">      �?   ħ �?[��<c�'>      �?   �k��?"���%>      �?   ���?݉@fR�8>      �?   ����?��T���:>      �?   T�!�?3&�F>      �?   � ��?<����[#>     ��?   �%�?�Y:/(A6>      �?   ����?��N��2>     ��?   8O�?�r�!'	>      �?   ��r�?���8{K>     ��?   �p��?9��l�9$>      �?   �
G�?�aj	�i9>     ��?   T|��?'\�|#<>      �?   $��?�}�dj�#>     ��?   �Wn�?׈MVx:>      �?   ,���?1�8o,>     ��?   D�$�?	c�/�
>      �?   @ |�?��x7|�1>     ��?   |���?��9>      �?   p #�?�IA��u=>     ��?   �s�?�x ٴ4>      �?   p���?edf�&�.>     ��?   ,�?��f���A>      �?   h�*�?v����2>     ��?   $gN�?RE\��K>      �?   �q�?'^��IE>     ��?   DΒ�?��&a��H>      �?   L���?�&KrQF>     ��?   ,���?�#/�'�>      �?   إ��?]X�c�?>     ��?    ��?�Ԯ}�>      �?   �e.�?�IdW�A>     ��?   �K�?���ΐ?>      �?   Xg�?��4*�A>     ��?   _��?�[�ǆJ>      �?   ���?1���0H>     ��?   ���?�hc#�]G>       @   ,*��?�Q�x
�F>     @ @   p���?ek�R�.N>     � @   �� �?�Ӿ�n@>     � @   �b�?�����O>      @   $Q/�?CJ���O>     @@   ��E�?������G>     �@   �[�?�3E�{A>     �@   T�p�?�SfI�S:>      @   X΅�?B6)�1�<>     @@   �3��?>ځ���7>     �@   $��?s(��N>     �@   @���?V�
6�f=>      @   (���?��{��>     @@   (W��?��-�Jg >     �@   ����?��"a�PK>     �@   xm�?,S��ڤ6>      @   ���?�6��hb">     @@    �-�?�k,�<>     �@   X�>�?�0����=>     �@   �O�?�׀IX�H>      @   �-_�?���
@>     @@   ��n�?���2E>     �@   �P~�?�=�ő�8>     �@   lj��?�[j&,>      @   L7��?��x��82>     @@   ����?c�#V�B>     �@   0��?7ڨ.�Y>     �@   P���?�[�p&>      @   ؔ��?h4�M��A>     @@   � ��?E�p�l E>     �@   �+��?�o�$�E>     �@   h��?\���*�K>      @   ���?-�?��B>     @@   P8�?�(l�|�@>     �@   �p!�?u���@�J>     �@   @p-�?�V��1>      	@   �89�?����5>     @	@   <�D�?��ƀ�7>     �	@   h)P�?R`D�OG>     �	@   �T[�?9%� ��K>      
@   �Mf�?��/�<>     @
@   �q�?�Ò��?>     �
@   �{�?4��2G<>     �
@   L��?Â���|/>      @   �Y��?���s�
@>     @@   �k��?��Ò�a@>     �@   XS��?x(3��u8>     �@   ���?v�O,ib>      @   ȥ��?�&L͒C>     @@   ���?��}��L>     �@   �X��?Lo����>     �@   �x��?-�Ϡ�9>      @   �s��?6FID?9>     @@   8J��?����gsL>     �@   d���?��y>     �@   ���?>�&�09C>      @   ����?
��<�A>     @@   (J�?I�V	C>     �@   `w�?��^@�N>     �@   ���?�#��%�@>      @   �s�? �M�K>     @@    D'�?ή�Q��->     �@   ��.�?9!���G>     �@   ��6�?.����1>      @   >�?.1�NcB>      @   �cE�?�sǔ�1>     @@   L�L�?�n�HN>     `@   H�S�?�W��$>     �@   8�Z�?
Ȃ�q�;>     �@   ��a�?N�/�[7>     �@   (�h�?�=�mC>     �@   0oo�?�H75M>      @   Hv�?P��.�#>      @   �|�?�G���7>     @@   �*��?�#4��2I>     `@   ����?o���oJ>     �@   ����?���-��#>     �@   ���?�h��%F>     �@   @��?R�x^D>     �@   PP��?�� s�@>      @   4L��?P�_!
�#>      @   4��?��:#�G>     @@   L��?qg�:&J>     `@   Hɹ�?5L$.��4>     �@   \w��?!�1�C>     �@   ���?���[<>     �@   D���?��<���=     �@   ���?��
~���=      @   �y��?������B>      @   ����?�~.���4>     @@   h��?��u�|�8>     `@   �E��?A8yL;>     �@   �h��?��41��C>     �@   �{��?-���+oF>     �@   $��?x���O>     �@   s��?�՝m�T2>      @   �W��?����=>      @   �-�?î�\�=>     @@   ��?���\=�=     `@   ��?j\&">     �@   �X�?��1�D>>     �@   ���?�#O#`�I>     �@   ��?�}���0>     �@   ��?���F\IE>      @   t{#�?��ׯ,B>      @   0�'�?�E� ]�$>     @@   ,>,�?��ކ?5>     `@   ��0�?��iIqE>     �@   ��4�?�ha�;>     �@   �9�?��A���D>     �@   �.=�?̤KF�w�=     �@   DMA�?�����=      @   `E�?ap�I0�H>      @   �gI�?��:���->     @@   �cM�?��%Q>     `@   @UQ�?Ly5ښoE>     �@   �;U�?v�g�0�/>     �@   �Y�?jv�U�G>     �@   �\�?�����yK>     �@   ,�`�?A%My��>      @   md�?���H>      @    h�?�p���M>     @@   0�k�?k��}<>     `@   �ho�?����f7O>     �@   ��r�?���}�O>     �@    �v�?+��i�I>     �@   @z�?�b�B'=>>     �@   `�}�?Z����M>      @   ����?1�����M>      @   �a��?R�~���=     @@   t���?QNT	��B>     `@   x��?�W3c�L>     �@   g��?�+(����=     �@   D���?q���J�K>     �@   L��?� ;,*>     �@   8!��?������D>      @   ,O��?� ����E>      @   Du��?��in]D>     @@   ����?%����3F>     `@   P���?^��F"VM>     �@   ����?�}�30}->     �@   @���?�~F	y�;>     �@   ����?l	R(>     �@   躰�?��\�7`>      @    ���?�dg���;>      @   ���?�;Sv�@E>     @@   <|��?�����M>     `@   �Y��?|}�;�2>     �@   ,0��?�<v��G>     �@   $ ��?̯�/p�">     �@   ����?���\(0>     �@   |���?[s$���F>      @   I��?�d�ӔV>      @   T���?���0)LK>     @@   h���?�)�5G�5>     `@   XY��?�|��zJ>     �@   @���?W�޾�L?>     �@   0���?����6:>     �@   <3��?��Q���B>     �@   x���?7o��/�M>      @   �Q��?�Kc�Z�0>      @   ����?�z-�A5>     @@   Z��?"B�DcI>     `@   ����?��`I�.>     �@    L��?L�d�%>     �@   ���?"�l"w �=     �@   �(��?�?��!>     �@   ���?��j^�J>      @   8���? ϞH��0>      @   LL��?���%�C>     @@   T���?��J�+N>     `@   d���?;l�>�0>     �@   �B��?�^{v�@>     �@   Ȋ��?�@Y˕B>     �@   @� �?T�l���0>     �@   ��?w4n4>      @    G�?�oN�=�;>      @   h|�?�L�{�/>     @@   <�	�?B�nu5>     `@   ���?���`�,+>     �@   d�?����5>     �@   �$�?l��  >     �@   �C�?~+^��M>     �@   �^�?�PK�QD >      @   ,u�?^{�#tF>      @   |��?�^4K�� >     @@   ���?��4�O
>>     `@   ���?XEړ� J>     �@   ���?(�gԹ�,>     �@   �� �?43-spF>     �@   ��"�?P`E5�+*>     �@   ��$�?=�QQ�D>       @-DT�!�?\3&��<e+000     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          �      	   m s c o r e e . d l l   CorExitProcess  k e r n e l 3 2 . d l l     FlsAlloc    FlsFree FlsGetValue FlsSetValue InitializeCriticalSectionEx CreateEventExW  CreateSemaphoreExW  SetThreadStackGuarantee CreateThreadpoolTimer   SetThreadpoolTimer  WaitForThreadpoolTimerCallbacks CloseThreadpoolTimer    CreateThreadpoolWait    SetThreadpoolWait   CloseThreadpoolWait FlushProcessWriteBuffers    FreeLibraryWhenCallbackReturns  GetCurrentProcessorNumber   GetLogicalProcessorInformation  CreateSymbolicLinkW SetDefaultDllDirectories    EnumSystemLocalesEx CompareStringEx GetDateFormatEx GetLocaleInfoEx GetTimeFormatEx GetUserDefaultLocaleName    IsValidLocaleName   LCMapStringEx   GetCurrentPackageId GetTickCount64  GetFileInformationByHandleExW   SetFileInformationByHandleW    0�   ��	   �
   @�   ��   �   @�   ��   �   P�   ��   �   ��   ̦   �    ا!   @�"   0�x   ��y   ��z   Ԫ�   ��   ��R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
         R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
         R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 4  
 -   i n c o n s i s t e n t   o n e x i t   b e g i n - e n d   v a r i a b l e s  
     D O M A I N   e r r o r  
     S I N G   e r r o r  
     T L O S S   e r r o r  
    
     r u n t i m e   e r r o r       R u n t i m e   E r r o r ! 
 
 P r o g r a m :     < p r o g r a m   n a m e   u n k n o w n >     . . .   
 
         M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y         atan2        �H��%%%��%��������HH����   p�   x�   ��   ��   ��   ��   ��   ��	   ��
   ��   Ⱥ   к   غ   �   �   �   ��    �   �   �   �    �   (�   0�   8�   @�   H�   P�   X�   `�    h�!   p�"   x�#   ��$   ��%   ��&   ��'   ��)   ��*   ��+   ��,   ��-   Ȼ/   л6   ػ7   �8   �9   �>   ��?    �@   �A   �C   �D    �F   (�G   0�I   8�J   @�K   H�N   P�O   X�P   `�V   h�W   p�Z   x�e   ��   ��  ��  ��  ��  ��  ��  ȼ  Լ  �	  �  ��  �  �  �  (�  4�  @�  L�  X�  d�  p�  |�  ��  ��  ��  ��  ��  Ľ  н  ܽ   �!  ��"   �#  �$  �%  $�&  0�'  <�)  H�*  T�+  `�,  l�-  ��/  ��2  ��4  ��5  ��6  ��7  ̾8  ؾ9  �:  �;  ��>  �?  �@   �A  ,�C  8�D  P�E  \�F  h�G  t�I  ��J  ��K  ��L  ��N  ��O  ��P  ȿR  ԿV  �W  �Z  ��e  �k  �l  ,��  8�  D�  P�  \�	  h�
  t�  ��  ��  ��  ��  ��  ��  ��,  ��;  ��>  �C  �k  (�  8�  D�  P�	  \�
  h�  t�  ��;  ��k  ��  ��  ��  ��	  ��
  ��  ��  ��;  �  �  $�  0�	  <�
  H�  T�  `�;  x�  ��	  ��
  ��  ��  ��;  ��  ��	  ��
  ��  �;  �   ,�	   8�
   D�;   P�$  `�	$  l�
$  x�;$  ��(  ��	(  ��
(  ��,  ��	,  ��
,  ��0  ��	0  ��
0  ��4   �	4  �
4  �8  $�
8  0�<  <�
<  H�@  T�
@  `�
D  l�
H  x�
L  ��
P  ��|  ��|  ����B   ػ,   ��q   p�    ���   ���   ���   ���   ���   ���   ��   ��    ��   ,��   8��   D��   P�C   \��   h��   t��   ��)   ���   ��k   ��!   ��c   x�   ��D   ��}   ���   ��   ��E   ��   ��G   ��   ��   �H   ��   ��   (��   4�I   @��   L��   ��A   X��   ��   h�J   ��   t��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��K   ���   ��   ��	   ��   ��   (��   4��   @��   L��   X��   d��   p��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��#   ��e   Ȼ*    �l   ��&   �h   Ⱥ
   �L   �.   $�s   к   0��   <��   H��   T�M   `��   l��   h�>   x��   0�7   ��   غ   ��N   �/   ��t   8�   ���   ��Z   �   ��O   ��(   ��j   p�   ��a   �   ��P   �   ���   ��Q   ��   �R   �-   �r    �1    �x   H�:   ,��    �   p�?   8��   H�S   �2   T�y   ��%   `�g   ��$   l�f   x��   л+   ��m   ���   `�=   ���   P�;   ���   ��0   ���   ��w   ��u   ��U   �   ���   ��T   ���   �   ��   (�6   �~   �    �V    �   ,�W   8��   D��   T��   d��   (�   t�X   0�   ��Y   X�<   ���   ���   ��v   ���   @�   ��[   ��"   ��d   ���   ���   ���   ��   ��   $��   H�   4�\   ���   @��   X��   p��   ���   P�   ���   ��]   �3   ��z   x�@   ���   8�8   ���   @�9   ���   X�   ��^   ��n   `�   �_    �5   �|   x�    �b   h�   (�`   �4   4��   L�{   ��'   d�i   p�o   |�   ���   ���   ���   ���   ���   ��F   ��p   a r     b g     c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     u k     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k   s y r   d i v       a r - S A   b g - B G   c a - E S   z h - T W   c s - C Z   d a - D K   d e - D E   e l - G R   e n - U S   f i - F I   f r - F R   h e - I L   h u - H U   i s - I S   i t - I T   j a - J P   k o - K R   n l - N L   n b - N O   p l - P L   p t - B R   r o - R O   r u - R U   h r - H R   s k - S K   s q - A L   s v - S E   t h - T H   t r - T R   u r - P K   i d - I D   u k - U A   b e - B Y   s l - S I   e t - E E   l v - L V   l t - L T   f a - I R   v i - V N   h y - A M   a z - A Z - L a t n     e u - E S   m k - M K   t n - Z A   x h - Z A   z u - Z A   a f - Z A   k a - G E   f o - F O   h i - I N   m t - M T   s e - N O   m s - M Y   k k - K Z   k y - K G   s w - K E   u z - U Z - L a t n     t t - R U   b n - I N   p a - I N   g u - I N   t a - I N   t e - I N   k n - I N   m l - I N   m r - I N   s a - I N   m n - M N   c y - G B   g l - E S   k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A   m i - N Z   a r - I Q   z h - C N   d e - C H   e n - G B   e s - M X   f r - B E   i t - C H   n l - B E   n n - N O   p t - P T   s r - S P - L a t n     s v - F I   a z - A Z - C y r l     s e - S E   m s - B N   u z - U Z - C y r l     q u z - E C     a r - E G   z h - H K   d e - A T   e n - A U   e s - E S   f r - C A   s r - S P - C y r l     s e - F I   q u z - P E     a r - L Y   z h - S G   d e - L U   e n - C A   e s - G T   f r - C H   h r - B A   s m j - N O     a r - D Z   z h - M O   d e - L I   e n - N Z   e s - C R   f r - L U   b s - B A - L a t n     s m j - S E     a r - M A   e n - I E   e s - P A   f r - M C   s r - B A - L a t n     s m a - N O     a r - T N   e n - Z A   e s - D O   s r - B A - C y r l     s m a - S E     a r - O M   e n - J M   e s - V E   s m s - F I     a r - Y E   e n - C B   e s - C O   s m n - F I     a r - S Y   e n - B Z   e s - P E   a r - J O   e n - T T   e s - A R   a r - L B   e n - Z W   e s - E C   a r - K W   e n - P H   e s - C L   a r - A E   e s - U Y   a r - B H   e s - P Y   a r - Q A   e s - B O   e s - S V   e s - H N   e s - N I   e s - P R   z h - C H T     s r     a f - z a   a r - a e   a r - b h   a r - d z   a r - e g   a r - i q   a r - j o   a r - k w   a r - l b   a r - l y   a r - m a   a r - o m   a r - q a   a r - s a   a r - s y   a r - t n   a r - y e   a z - a z - c y r l     a z - a z - l a t n     b e - b y   b g - b g   b n - i n   b s - b a - l a t n     c a - e s   c s - c z   c y - g b   d a - d k   d e - a t   d e - c h   d e - d e   d e - l i   d e - l u   d i v - m v     e l - g r   e n - a u   e n - b z   e n - c a   e n - c b   e n - g b   e n - i e   e n - j m   e n - n z   e n - p h   e n - t t   e n - u s   e n - z a   e n - z w   e s - a r   e s - b o   e s - c l   e s - c o   e s - c r   e s - d o   e s - e c   e s - e s   e s - g t   e s - h n   e s - m x   e s - n i   e s - p a   e s - p e   e s - p r   e s - p y   e s - s v   e s - u y   e s - v e   e t - e e   e u - e s   f a - i r   f i - f i   f o - f o   f r - b e   f r - c a   f r - c h   f r - f r   f r - l u   f r - m c   g l - e s   g u - i n   h e - i l   h i - i n   h r - b a   h r - h r   h u - h u   h y - a m   i d - i d   i s - i s   i t - c h   i t - i t   j a - j p   k a - g e   k k - k z   k n - i n   k o k - i n     k o - k r   k y - k g   l t - l t   l v - l v   m i - n z   m k - m k   m l - i n   m n - m n   m r - i n   m s - b n   m s - m y   m t - m t   n b - n o   n l - b e   n l - n l   n n - n o   n s - z a   p a - i n   p l - p l   p t - b r   p t - p t   q u z - b o     q u z - e c     q u z - p e     r o - r o   r u - r u   s a - i n   s e - f i   s e - n o   s e - s e   s k - s k   s l - s i   s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l   s r - b a - c y r l     s r - b a - l a t n     s r - s p - c y r l     s r - s p - l a t n     s v - f i   s v - s e   s w - k e   s y r - s y     t a - i n   t e - i n   t h - t h   t n - z a   t r - t r   t t - r u   u k - u a   u r - p k   u z - u z - c y r l     u z - u z - l a t n     v i - v n   x h - z a   z h - c h s     z h - c h t     z h - c n   z h - h k   z h - m o   z h - s g   z h - t w   z u - z a       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       @�P�L���Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy HH:mm:ss    S u n   M o n   T u e   W e d   T h u   F r i   S a t   S u n d a y     M o n d a y     T u e s d a y   W e d n e s d a y   T h u r s d a y     F r i d a y     S a t u r d a y     J a n   F e b   M a r   A p r   M a y   J u n   J u l   A u g   S e p   O c t   N o v   D e c   J a n u a r y   F e b r u a r y     M a r c h   A p r i l   J u n e     J u l y     A u g u s t     S e p t e m b e r   O c t o b e r   N o v e m b e r     D e c e m b e r     A M     P M     M M / d d / y y     d d d d ,   M M M M   d d ,   y y y y   H H : m m : s s                       8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7      �?5�h!���>@�������             ��      �@      �                          �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC                                            �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               �       �      ��      ������    ����    ��      ��            8C      8C      0<      0<��+eGW@��+eGW@  ��B.�?  ��B.�?:;����=:;����=�ѱt�?Z�fUUU�?���&WU�?{������?                Mu�{�<`�w>�,  �g5RҌ<t�ӰY  a��aN�`<țuE�  l{�]���<��lX�  ќ/p=�><���2��  ؼcnQ�<P[� {8�&TŤ<�-���B �?RbSQ�<zQ}<�r �S?���<u�o�[� _/:>��<��h1�� �æDAo�<֌b�; �������<8bunz8 ���+G�<�|�eEk 1�	m���<����� �
r�7�<䦅� ���MuM�<�1
� J��]9ݏ<�d�< )}̌/�<ʩ:7�q �^�s)ҧ<���4ۧ mL*�H��<"4L�� ��%F��<).�!
 ��`�cC<-�a`N y����n<�<���� ��z�ΐv<'*6�ڿ 	*(�̃�<�,�v�� ���	�<�O�V+4 ���5�<�'�6Go 	T��c�<)TH�� 5�d+�2�<H!�o� 
���<�U:�~$ �s ��<$"U�8b qU�M��<�;f�� �GΆ�+�<.e<�� �o � �<s_��u ���"a�<�gBV�_ ��F�D�<��s� Ul֫��e<bN�6�� �g�����<�L��% ���<�D��h ����/��<۠*B� D_�Y��{<6w��� <(��`�<��Ͱ77	 �b� ��<ONޟ�}	 'Α+��q<�𣂑�	 �.�X4m�<d�]{f
 ����|'�<\%>�U
 �Zsn�i�<��yUk�
 �3˒w�<��Z���
 �-�f$�<�O��3 ���.�<F^��v ��_
��t<��K�� ��0�ns<�R�ݛ �Y	я��<K�W.�g h�l,kg<i��� � ���6	p�<{�J- �=���t<����X ����PZ�<�2�� ��Js��<^�{3�� ӈ:`�t<�?��.P &I	�'o�<ِ����  �A�Î<'Za�� ��1�d�<@En[vP �͑M;�w<ؐ����       �?       �9��B.�@  ׽2b      �        �������         0<  0<�dW�dW       ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          A6]�b�q7            �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �sinh    cosh    tanh    atan2   fabs    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter  \<h<p<|<�<�<�<�<�<�<�<�<�<���<�< ========(=,=0=4=��8=<=@=D=0�H=L=P=T=X=\=�`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=><>\>|>�>�>�> ? ?H?d?t?x?�?�?�?�?�?�?�?@<@d@�@�@�@�@AHAtA���A�A�A�A�A__based(    __cdecl __pascal    __stdcall   __thiscall  __fastcall  __vectorcall    __clrcall   __eabi  __ptr64 __restrict  __unaligned restrict(    new     delete =   >>  <<  !   ==  !=  []  operator    ->  *   ++  --  +   &   ->* /   <   <=  >   >=  ,   ()  ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall' `typeof'    `local static guard'    `string'    `vbase destructor'  `vector deleting destructor'    `default constructor closure'   `scalar deleting destructor'    `vector constructor iterator'   `vector destructor iterator'    `vector vbase constructor iterator' `virtual displacement map'  `eh vector constructor iterator'    `eh vector destructor iterator' `eh vector vbase constructor iterator'  `copy constructor closure'  `udt returning' `EH `RTTI   `local vftable' `local vftable constructor closure'  new[]   delete[]   `omni callsig'  `placement delete closure'  `placement delete[] closure'    `managed vector constructor iterator'   `managed vector destructor iterator'    `eh vector copy constructor iterator'   `eh vector vbase copy constructor iterator' `dynamic initializer for '  `dynamic atexit destructor for '    `vector copy constructor iterator'  `vector vbase copy constructor iterator'    `managed vector copy constructor iterator'  `local static thread guard'  Type Descriptor'    Base Class Descriptor at (  Base Class Array'   Class Hierarchy Descriptor'     Complete Object Locator'   U S E R 3 2 . D L L     MessageBoxW GetActiveWindow GetLastActivePopup  GetUserObjectInformationW   GetProcessWindowStation           8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �        ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               ( ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                                                            �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#SNAN  1#IND   1#INF   1#QNAN  C O N O U T $   A      H                                                           � �   RSDSxwnڤ)E�'�'ҔN�   E:\repos\cmNodes\src\obj\cmnodes_r14_Win32_Release.pdb      �   �                      �l�lm    X�       ����    @   �lp�        ����    @   0m           @mm               Xmdmm    ��       ����    @   Hm            ���m           �m�mm    ��       ����    @   �m           �m�m�lm    ��       ����    @   �m           n(n�lm    ��       ����    @   n��       ����    @   `n           pnDn�n�n    �       ����    @   �n           �n�n�n    ,�        ����    @   �n           �n�n                D� o           oo8o    D�       ����    @    o`�        ����    @   To           do8o                |��o           �o�oDn�n�n    |�       ����    @   �o            ���o           �o�odmm    ��       ����    @   �o            ��$p           4pHpdp�lm    ��       ����    @   $p��       ����    @   �p           �pdp�lm                ���p           �p�pdp�lm    ��       ����    @   �p            �q           q(q�lm    �       ����    @   q            (�Xq           hq|q�m�lm    (�       ����    @   Xq            D��q           �q�q�q�lm    D�       ����    @   �q`�       ����    @   r           r�q�lm                |�<r           Lr`r�q�lm    |�       ����    @   <r            ���r           �r�r�q�lm    ��       ����    @   �r            ���r           �rs�q�lm    ��       ����    @   �r            ��8s           Hs\s�q�lm    ��       ����    @   8s            ���s           �s�s�q�lm    ��       ����    @   �s            ��s           �st�q�lm    �       ����    @   �s            (�4t           DtXt�q�lm    (�       ����    @   4t            D��t           �t�t�q�lm    D�       ����    @   �t            `��t           �t u�q�lm    `�       ����    @   �t            |�0u           @uTu�q�lm    |�       ����    @   0u            ���u           �u�u�q�lm    ��       ����    @   �u            ���u           �u�u�q�lm    ��       ����    @   �u            ��,v           <vPv�q�lm    ��       ����    @   ,v            ���v           �v�v�q�lm    ��       ����    @   �v            ��v           �v�v�q�lm    �       ����    @   �v            0�(w           8wLw�q�lm    0�       ����    @   (w            L�|w           �w�w�q�lm    L�       ����    @   |w            h��w           �w�w�q�lm    h�       ����    @   �w            ��$x           4xHx�q�lm    ��       ����    @   $x            ��xx           �x�x�q�lm    ��       ����    @   xx            ���x           �x�x�q�lm    ��       ����    @   �x            �� y           0yDy�q�lm    ��       ����    @    y            ��ty           �y�y�q�lm    ��       ����    @   ty            ��y           �y�y�q�lm    �       ����    @   �y            8�z           ,z@z�q�lm    8�       ����    @   z            X�pz           �z�z�q�lm    X�       ����    @   pz            t��z           �z�z�q�lm    t�       ����    @   �z            ��{           ({<{�q�lm    ��       ����    @   {            ��l{           |{�{�q�lm    ��       ����    @   l{            ���{           �{�{�q�lm    ��       ����    @   �{            ��|           $|8|�q�lm    ��       ����    @   |            �h|           x|�|�q�lm    �       ����    @   h|             ��|           �|�|�q�lm     �       ����    @   �|            @�}            }4}�q�lm    @�       ����    @   }            `�d}           t}�}�q�lm    `�       ����    @   d}            ���}           �}�}�q�lm    ��       ����    @   �}            ��~           ~,~�mm    ��       ����    @   ~            ��\~           l~|~�mm    ��       ����    @   \~            ���~           �~�~�mm    ��       ����    @   �~             ��~           �mm     �       ����    @   �~             �L           \l�mm     �       ����    @   L            D��           ���mm    D�       ����    @   �            h��           ���mm    h�       ����    @   �            ��<�           L�\��mm    ��       ����    @   <�            ����           �����mm    ��       ����    @   ��            ��܀           ����mm    ��       ����    @   ܀            ��,�           <�L��mm    ��       ����    @   ,�            �|�           �����mm    �       ����    @   |�            <�́           ܁��mm    <�       ����    @   ́            \��           ,�<��mm    \�       ����    @   �            |�l�           |����mm    |�       ����    @   l�            ����           ̂܂�mm    ��       ����    @   ��            ���           �,��mm    ��       ����    @   �            ��\�           l�|��mm    ��       ����    @   \�            ���           ��̃�mm    �       ����    @   ��            @���           ���mm    @�       ����    @   ��            h�L�           \�l��mm    h�       ����    @   L�            ����           �����mm    ��       ����    @   ��            ���           ����mm    ��       ����    @   �            ��<�           L�\��mm    ��       ����    @   <�            ���           �����mm    �       ����    @   ��            @�܅           ����mm    @�       ����    @   ܅            h�,�           <�L��mm    h�       ����    @   ,�            ��|�           �����mm    ��       ����    @   |�            ��̆           ܆��mm    ��       ����    @   ̆            ���           ,�<��mm    ��       ����    @   �            �l�           |����mm    �       ����    @   l�            <���           ̇܇�mm    <�       ����    @   ��            l��           �,��mm    l�       ����    @   �            ��\�           l�|��mm    ��       ����    @   \�            ����           ��̈�mm    ��       ����    @   ��            ����           ���mm    ��       ����    @   ��            �L�           \�l��mm    �       ����    @   L�            H���           �����mm    H�       ����    @   ��            t��           ����mm    t�       ����    @   �            ��<�           L�\��mm    ��       ����    @   <�            ����           �����mm    ��       ����    @   ��            ��܊           ����mm    ��       ����    @   ܊             �,�           <�L��mm     �       ����    @   ,�            L�|�           �����mm    L�       ����    @   |�            x�̋           ܋��mm    x�       ����    @   ̋            ���           ,�<��mm    ��       ����    @   �            ��l�           |����mm    ��       ����    @   l�            ���           ̌܌�mm    �       ����    @   ��            ,��           �,��mm    ,�       ����    @   �            X�\�           l�|��mm    X�       ����    @   \�            ����           ��̍�mm    ��       ����    @   ��            ����           ���mm    ��       ����    @   ��            ��L�           \�l��mm    ��       ����    @   L�            ���           �����mm    �       ����    @   ��            0��           ����mm    0�       ����    @   �           8�H��mm    X�       ����    @   (�            ��x�           ����H��mm    ��       ����    @   x�            ��̏           ܏��H��mm    ��       ����    @   ̏            �� �           0�D�H��mm    ��       ����    @    �            �t�           ����H��mm    �       ����    @   t�            4�Ȑ           ؐ�H��mm    4�       ����    @   Ȑ            `��           ,�@�H��mm    `�       ����    @   �            ��p�           ����H��mm    ��       ����    @   p�            ��đ           ԑ�H��mm    ��       ����    @   đ            ���           (�<�H��mm    ��       ����    @   �            �l�           |���H��mm    �       ����    @   l�            <���           Вܒ8o    <�       ����    @   ��            `��           �(��n    `�       ����    @   �            ��X�           h�x��mm    ��       ����    @   X�            ����           ��ē�n    ��       ����    @   ��            ����           ���mm    ��       ����    @   ��            ��D�           T�`�|�    ��       ����    @   D��        ����    @   ��           ��|�                ,�Ĕ           Ԕ�(n�lm    ,�       ����    @   Ĕ            `�r            p�0m            ���            ��n            ,��n            `�To            H���           �����n    H�       ����    @   ��            ��`n            d��            ��    d�        ����    @   �            |�8�           H�P�    |�        ����    @   8�            ����           ����P�    ��       ����    @   ��            ���p            ����           ���    ��        ����    @   ��            �  �R 0y                     ����    ����    ����    s�    ����    ����    �����%�    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    '�����    3�����    ����    ����    ������    ������    ����    ����    �    ����    |���    ����    ��    ����    ����    ����    �
    ����    ����    ����        ����    ����    ����    y    ����    ����    ����    h    ����    ����    ����         ����    ����    ����    �!    ����    ����    �����O�O    ����    ����    ����    �Q    ����    ����    ����y\�\    ����    ����    ����]]    ����    ����    ����    =k    ����    ����    ����    �l        �l����    ����    ����    bm    ����    ����    ����    A{    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    {�                ��DT    ��          �� �� �� R    cmnodes_r14.cdl c4d_main  ��         R�  �                     � �� � � 4� D� P� \� x� �� �� �� �� Ҝ � �� �  � .� F� X� n� �� �� �� ҝ � � &� N� V� j� ~� �� �� �� �� Ğ О � � � � 2� B� T� h� z� �� �� �� �� �� ̟ ڟ �  � � "� 6� D�     !EncodePointer � DecodePointer �GetCommandLineA GetCurrentThreadId  PGetLastError  3HeapFree  /HeapAlloc mIsProcessorFeaturePresent gIsDebuggerPresent 
SetLastError  QExitProcess fGetModuleHandleExW  �GetProcAddress  �MultiByteToWideChar �WideCharToMultiByte �GetProcessHeap  �GetStdHandle  >GetFileType DeleteCriticalSection �GetStartupInfoW bGetModuleFileNameA  -QueryPerformanceCounter 
GetCurrentProcessId �GetSystemTimeAsFileTime 'GetEnvironmentStringsW  �FreeEnvironmentStringsW �UnhandledExceptionFilter  ASetUnhandledExceptionFilter HInitializeCriticalSectionAndSpinCount PSleep 	GetCurrentProcess _TerminateProcess  qTlsAlloc  sTlsGetValue tTlsSetValue rTlsFree gGetModuleHandleW  �WriteFile cGetModuleFileNameW  8HeapSize  �LCMapStringW  %EnterCriticalSection  �LeaveCriticalSection  �GetConsoleCP  �GetConsoleMode  �SetFilePointerEx  rIsValidCodePage �GetACP  �GetOEMCP  �GetCPInfo ?RaiseException  �RtlUnwind �LoadLibraryExW  6HeapReAlloc �OutputDebugStringW   SetStdHandle  �WriteConsoleW �GetStringTypeW  �FlushFileBuffers  � CreateFileW  CloseHandle KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                 N�@���Du�  s�     ��                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                acos            atan            cos                   �?pow     sin             sqrt    ?  ?  �[�[�[�[�[�[�[�[�[�[����    �����
                                                          ����            asin            log     @�    @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                            0��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��               C   T�X�\�`�d�h�l�p�x����������������������������������������� ������ �,�4�@�L�P�T�`�t�       ������������������������� �4�<�D�L�T�\�d�l�t�|�������������T�����������0�D�L�T�h������                                   T�            T�            T�            T�            T�                          ؾ        pd�hxjX�                        �����&     d�   h�   X�   \�   `:   h:!   p:   l�   t�   ��   x:   ��   ��   ��    ��   ��   ��   �:   ��   �:   �:   �:   �:   �:"   �:#   �:$   �:%   �:&   �:      �      ���������              �       �D        � 0                                                                                                                                                                                                                                                                                           ؾ.   Ծ � � � � � � � � �(�$�$�$�$�$�$�$�.   pdrf             �            tf   ���5      @   �  �   ����             ����         �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                  �$c    .?AVNodeData@@  $c    .?AVBaseData@@  $c    .?AVCustomGuiData@@ $c    .?AVCommandData@@   $c    .?AVSceneHookData@@ $c    .?AVShaderData@@    $c    .?AViCustomGui@@    $c    .?AVSubDialog@@ $c    .?AVGeDialog@@  $c    .?AVcmMenuButton@@  $c    .?AVGeUserArea@@    $c    .?AVcmRealDlg@@ $c    .?AVcmRealGui@@ $c    .?AVcmPrefsObject@@ $c    .?AVPrefsDialogObject@@ $c    .?AVcmNodesPrefsObject@@    $c    .?AVcmNodeTree@@    $c    .?AVcmNodeForest@@  $c    .?AVcmNodeOutput@@  $c    .?AVcmNodeBase@@    $c    .?AVcmNodeMaterial@@    $c    .?AVcmNodeTexture@@ $c    .?AVcmNodeColor@@   $c    .?AVcmNodeShuffle@@ $c    .?AVcmNodeCopy@@    $c    .?AVcmNodeBlend@@   $c    .?AVcmNodeMath@@    $c    .?AVcmNodeClamp@@   $c    .?AVcmNodeCurves@@  $c    .?AVcmNodeGrade@@   $c    .?AVcmNodeColorspace@@  $c    .?AVcmNodeFilter@@  $c    .?AVcmNodeColorize@@    $c    .?AVcmNodeInvert@@  $c    .?AVcmNodeTransform@@   $c    .?AVcmNodeDistort@@ $c    .?AVcmNodeEmboss@@  $c    .?AVcmNodeMatrix@@  $c    .?AVcmNodeBlur@@    $c    .?AVcmNodeEdgeDetect@@  $c    .?AVcmNodeDirBlur@@ $c    .?AVcmNodeHighPass@@    $c    .?AVcmNodeInfo@@    $c    .?AVcmNodeSpecular@@    $c    .?AVcmNodeDistance@@    $c    .?AVcmNodeSwitch@@  $c    .?AVcmNodeReflection@@  $c    .?AVcmNodeNoop@@    $c    .?AVcmNodeDiffuse@@ $c    .?AVcmNodeFresnel@@ $c    .?AVcmNodeTiler@@   $c    .?AVcmNodeShadow@@  $c    .?AVcmNodeNormalMap@@   $c    .?AVcmNodeCondition@@   $c    .?AVcmNodeProjector@@   $c    .?AVcmNodeVrayAdvanced@@    $c    .?AVcmNodeCmd_Cut@@ $c    .?AVcmNodeCmd_Copy@@    $c    .?AVcmNodeCmd_Paste@@   $c    .?AVcmNodeCmd_Delete@@  $c    .?AVcmNodeCmd_SelectAll@@   $c    .?AVcmNodeCmd_DeselectAll@@ $c    .?AVcmNodeCmd_Disconnect@@  $c    .?AVcmNodeCmd_FrameSelected@@   $c    .?AVcmNodeCmd_Prefs@@   $c    .?AVcmNodeCmd_AddTree@@ $c    .?AVcmNodeCmd_TreeMenu@@    $c    .?AVcmNodeCmd_NodeMenu@@    $c    .?AVcmNodeCmd_ZoomIn@@  $c    .?AVcmNodeCmd_ZoomOut@@ $c    .?AVcmNodeCmd_Zoom100@@ $c    .?AVcmNodeCmd_ResetView@@   $c    .?AVcmNodeCmd_CalcPreview@@ $c    .?AVcmNodeCreateCmd_NodeSolidColor@@    $c    .?AVcmNodeCreateCmd_NodeTexture@@   $c    .?AVcmNodeCreateCmd_NodeClamp@@ $c    .?AVcmNodeCreateCmd_NodeColorspace@@    $c    .?AVcmNodeCreateCmd_NodeCurves@@    $c    .?AVcmNodeCreateCmd_NodeFilter@@    $c    .?AVcmNodeCreateCmd_NodeGrade@@ $c    .?AVcmNodeCreateCmd_NodeMath@@  $c    .?AVcmNodeCreateCmd_NodeBlend@@ $c    .?AVcmNodeCreateCmd_NodeCopy@@  $c    .?AVcmNodeCreateCmd_NodeShuffle@@   $c    .?AVcmNodeCreateCmd_NodeBlur@@  $c    .?AVcmNodeCreateCmd_NodeDirBlur@@   $c    .?AVcmNodeCreateCmd_NodeDistort@@   $c    .?AVcmNodeCreateCmd_NodeEdgeDetect@@    $c    .?AVcmNodeCreateCmd_NodeEmboss@@    $c    .?AVcmNodeCreateCmd_NodeMatrix@@    $c    .?AVcmNodeCreateCmd_NodeNormalMap@@ $c    .?AVcmNodeCreateCmd_NodeTransform@@ $c    .?AVcmNodeCreateCmd_NodeOutput@@    $c    .?AVcmNodeCreateCmd_NodeMaterial@@  $c    .?AVcmNodeCreateCmd_NodeColorize@@  $c    .?AVcmNodeCreateCmd_NodeInfo@@  $c    .?AVcmNodeCreateCmd_NodeHighPass@@  $c    .?AVcmNodeCreateCmd_NodeSwitch@@    $c    .?AVcmNodeCreateCmd_NodeInvert@@    $c    .?AVcmNodeCreateCmd_NodeSpecular@@  $c    .?AVcmNodeCreateCmd_NodeVrayAdvanced@@  $c    .?AVcmNodeCreateCmd_NodeDistance@@  $c    .?AVcmNodeCreateCmd_NodeReflection@@    $c    .?AVcmNodeCreateCmd_NodeNoop@@  $c    .?AVcmNodeCreateCmd_NodeDiffuse@@   $c    .?AVcmNodeCreateCmd_NodeFresnel@@   $c    .?AVcmNodeCreateCmd_NodeTiler@@ $c    .?AVcmNodeCreateCmd_NodeShadow@@    $c    .?AVcmNodeCreateCmd_NodeCondition@@ $c    .?AVcmNodeCreateCmd_NodeProjector@@ $c    .?AVcmNodeCreateCmd_NodeInput@@ $c    .?AVcmTreeBookmarkCmd_Bookmark@@    $c    .?AVcmTreeBookmarkCmd_Bookmark0@@   $c    .?AVcmTreeBookmarkCmd_Bookmark1@@   $c    .?AVcmTreeBookmarkCmd_Bookmark2@@   $c    .?AVcmTreeBookmarkCmd_Bookmark3@@   $c    .?AVcmTreeBookmarkCmd_Bookmark4@@   $c    .?AVcmTreeBookmarkCmd_Bookmark5@@   $c    .?AVcmTreeBookmarkCmd_Bookmark6@@   $c    .?AVcmTreeBookmarkCmd_Bookmark7@@   $c    .?AVcmTreeBookmarkCmd_Bookmark8@@   $c    .?AVcmTreeBookmarkCmd_Bookmark9@@   $c    .?AVcmNodeEditorUserArea@@  $c    .?AVcmNodeEditorDialog@@    $c    .?AVcmNodeEditorCommand@@   $c    .?AVcmTreeManagerDialog@@   $c    .?AVcmTreeManagerCommand@@  $c    .?AVcmUpdateNodeThread@@    $c    .?AVC4DThread@@ $c    .?AVcmNodeShader@@  $c    .?AVGeModalDialog@@ $c    .?AVNeighbor@@  $c    .?AVGeListView@@    $c    .?AVSimpleListView@@    $c    .?AVtype_info@@                                                                                                                                                                                                                                                                                                                    $  040T0a0}0�0�0�0�0�0�0�0�0�0�011*1>1W1h1y1�1�1�1�1�1�1�12"2.2<2P2i2�2�2�2�2�2�2�233&3:3S3p3�3�3�3�3�3�3�344$4=4Z4k4w4�4�4�4�4�4�4�45'5;5L5X5f5~5�5�5�5�566/6a6r6�6�6�6�6�6&7c7t7�7�7�7�7�78$888e8�8�8�8�8�8�8
99D9V9`9n9w9�9�9�9�9�9�9�9:-:A:f:p:�:/;c;�<�<�<�<�=�=�=�=>a>i>z>    �   0W0�01x1�12x2�23Q3�3�4�45�5�5�6�6G7w7�7?8@9H9�9�9�9�9�9 :�:�: ;;B;J;d;�;�;�;�;�;'<n<<�<�<==W=�=�=�=�=�=>>G?Z?b?�?�?�?�?   0  �   �0�0�011�1�1�12G2^2k2�3�304\4�7�78e8�8999{9�9�9�9i:w:�:�:�:�:�:�:�:�:;#;+;3;S;z;�;�;�;�;<F<`<�<�<�<4=I=Z=z=�=�=�=�=�=�=>a>�>�> ? ?�?�? @    �0�0�01131D1{1�2�2�2�2�283G3\3�3�3�3�3�3�3@4X4k4�4�4�455V5e5w5�5�5�5�5656M6�6�67$797p7}7�7�7�7�7�788Q8Y8�8�8�8/:C:K:S:y:�:�:�:�:�:�:�:;%;-;R;Z;~;�;�;�;�;�;�;�;<C<P<f<s<�<�<�<�<�<�<�<�<�<�<=!=2=Q=b=n=|=�=�=�=�=�=�=>4>J>S>s>�>�>�>�>�>�>�>?!?5?J?[?l?}?�?�?�?�?�?�?   P  |  0010B0T0t0�0�0�0�0�0�0�01131H1^1r1�1�1�1�1�1�1�122/2E2Y2n22�2�2�2�2�2�2
3353I3^3o3�3�3�3�3�344$4;4L4]4i4�4�4�4�4�4�4�455$505>5O5d5x5�5�5�5�5�566-6L6]6n66�6�6�6�6�6�6�67$7C7T7e7v7�7�7�7�7�7�7�78/8@8q8~8�8�8�8�8�8�8'9n99�9�9�9�9�9�9�9>:E:	;;6;P;i;�;�;�;�;�;<!<5<N<h<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======�=�=�=>7>O>b>�>�>�>�>�>?'???R?u?�?�?�?�?�?   `  h  0)0<0_0}0�0�0�0�011,1O1m1�1�1�1�1�12"2E2c2{2�2�2�2�2�2�23333H3i3~3�3�3�3�34&464K4c4x4�4�4�4�4�4�45535H5^5n5�5�5�5�5�5�566.6>6S6k67d7�7�7�7�7�7�7	88878=8b8�8�8�8�8�899"9D9J9g9�9�9�9�9�9:5:K:q:�:�:�:�:�:�:;";8;d;�;�;�;�;�;�;�;�;<#<,<K<m<v<�<�<�<�<�<�<�<==$=@=Q=`=v=�=�=�=�=�=�=>>!>->;>L>X>}>�>�>�>�>�>�>??%?3?D?P?u?�?�?�?�?�?�?�? p  �   00"0>0c0l0}0�0�0�0�0�0�0�01161G1V1l1}1�1�1�1�1�1�1�1k4�4�45[5�5�5�5�5�56 6(6=6S6_6s6�6�6�67d7�7�7�7�788T8�8�8�8E9\9t9�9�9�:�:�:!;�;�;�;�;�;�; <<'<9<J<[<p<�<�<�<�<�<==(=;=G=s=�=�=�=�=�=>>>W>h>y>�>�>�>�>??-?9?^?o?�?�?�?�?�?   �  l  0,060D0J0b0h0�0�0�0�0�0�0�0�0�0
1"1(1@1U1�1�1�1�1�1�122/2@2Z2k22�2�2�2�2�2�23$353P3m3�3�3�3�3�3�3 4474H4a44�4�4�4�4�45 595W5h5�5�5�5�5�5�56/6@6Y6w6�6�6�6�6�67717O7`7y7�7�7�7�7�7	8'888Q8o8�8�8�8�8�8�89)9G9X9q9�9�9�9�9�9::0:I:g:x:�:�:�:�:�:;!;?;P;i;�;�;�;�;�;�;<(<A<_<p<�<�<�<�<�< ==7=H=a==�=�=�=�=�=>:>I>X>�>�>�>�>�>??%?e?v?�?�?�?�?�?�? �  �   0070A0Y0s0�0�0�0�0�0�011<1P1a1�1�12%2D2U2�2�2�2�2F3Z3�3�3�3�34-464R5Z5h5�5�5�5�5�5�5�5�566L6\6�6�6�67N7]7q7�7�7�7�7�7�7�78!8,848j9v9�9�9�<==*=�=>>H>x>�>�>?H?x?�?�?   �  �   080h0�0�0X1�1�1�1�12H2x2�2�2383h3�3�3�3(4X4�4�45H5x5�5�5�5(6X6�6�6+7h7�7�7�7�7'8G8`8q8}8�8�8�89D9h9p9�9�9�9�9:):T:a:�:�:�:�:$;F;d;�;�;�;$<H<P<t<�<�<�<==%=T=x=�=�=�=�=�=> >D>g>s>�>�>�>?4?X?`?�?�?�?   �  �   0(000T0v0�0�0�0�0141U1]1�1�1�1�122D2c2s2�2�2�2333T3x3�3�3�34'434t4�4�4�4�4545Y5o5z5�5�5�5�56#646S6h6�6�6�67787�7�7�78�8�8�8�8Y;j;|;�;?<P<\<x<�<�<�<�<�<�<�< =1=B=N=o=�=�=�=�=�=�=�=>#>4>@>a>r>�>�>�>�>�>�>�>?!?-?N?i?z?�?�?�?�?�?   �  �    0�0D1H1L1P1T1X1\1`1d1h1l1p1t1x1�1�1�1�1�1�1�1�1 2222222.2�2�2�2�2�2�2�2�2�2�2�2�2�2�23/3Q3r3�3�34x5�578g8�9:�:�:�:�:;";C;X;�; <"<P<x<�<�<?�?   �  �   �0�0�0�12=2|2�2�2�2�2�2 3<3X3t3�34�4�4�4�4G5l5�566@6Q6�67#7I7Z7�7�7	88V8^8l88�8�899�9�9�9�9:}:�:�:�:�:�:�:�:�:�:�:;;%;3;\;m;y;�;�;�;�;�;<<"<0<E=i=�=�=�=>">.><>X>g>�>�>�>�>�>�>?6?M?o?�?�?�?�?   �    0G0[0�01(1o1�1�1�1�1�1�122(262G2�2�2�23-3U3o3�3�3�34:4[4}4�4�4�455&5T5w5�5�5�5�5�5686�6�6�6�6%7?7�7�7�7�78(898h8�9�9::�:�:�:�:�:;;';k;�;�;<<<h<y<�<�<�<�<#=�=�=�=�=�=�=�=�=�=�=X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �  �   0&0/0N0_0p0|0�0K1\1h1�1�1�1�12S2d2p2�2333=3N3_3k3�3"4]4x4�4�4�4�4�4�45%515?5k5|5�5�5�5�5�5�5Q6q6�6�6�6=7]7�7�7�7818M8n8�8�8�8D9S9q9�9�9.:o:�:�:	;5;w;�;�;�;<j<�<�<1=w=�=�=�=�=�=>>7>g>x>�>�>�>�>�>�> ??�?�?�?�?     H   0U0f0r0�0�0�0�0�0�031�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5#5*5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5<6�677 7�7�7�7�78�8�8�8�859F9R9`9�9:A:[:�;3<�<�<8=X=�=#>B>�>�>�>??\?d?�?�?�?    p   :0�0K1�1�1,343�6�67'7�7�7C8s8�89909F9Z9�9�9:�:;-;z;�;�;�;�;�;�;�<i=�=�=�=5>l>�>�>�>�>??R?^?o?�?�?   �   11g1o1w11�1�1=2u2�2�2�233�3p4�4�4�4�4 535E5�5�5�5�5�5�6�6�6767�7�7�7�78(8s8�8"9d9::L:�:�:�:�:�:�:;>;�;�;�;�;�;�;�<�<�<�<@=d=r=~=�=�=>$>�>�>2?�?�?�?�?   0 P   I0r0�01�1�12!2�2�23�3	4L4T4�4�5�5�5�5�617a7n7�7�7�7�9s:;|;�;�;s<�<�< @ �   B4a4�4�455&575C5�5�5�5�5�5E6V6b6p6�6�6�6�6�6	77�7�7�7�7�8�8�9�9d:y:�:�:�:�:�:�:�: ;;;+;=;Z;k;w;�;�;�;�;�;�;�;<<<<!<�<�<�=(>8>_>u>�>�>C?]?�?�?   P �   +0E0�0�01-1�1�1�12o2�2�2�2W3q3�3�3?4Y4�4�4&5_5�5�5676T6�6�67�7�7�7%8s8�8�8%9[9`9~9�9�9�9:4:t:x:|:�:�:�:;B;l;�;<Q<e<w<�<�<�<�<�<�<={=�=>+>>�>�>�>�>?5?D?Y?y?�?�?�?�?   ` �   0_0u0�0�0�0�01$191Y1�1�1�1�1�192D23B3J3�3�3�34�4�445W5]5z5�5�5�5�56(6E6b66�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6,70747T8x8~8�8�8929_9�9�9�9:@:m:�:�:�:!;N;{;�;�;</<\<�<�<�<===j=�=�=�=>K>x>�>�>�>,?Y?�?�?�?   p �  0:0g0�0�0�01H1u1�1�1�1)2V2�2�2�2
373d3�3�3�34E4o4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666666636D6P6y6�6�6�6�6#757<7N7T77�7�7�7�7�768H8O8a8h8z8�8�8�8�8�8�869H9O9a9h9z9�9�9�9�9�9::0:G:^:u:�:�:�:�:�:�:�:�:�:�:�:�:�:;;';m;|;�;�;�;�;�;�;<<)<:<L<_<w<�<�<===5=I=[=l=}=�=�=�=�=>>4>K>b>y>�>�>�>�>�>??1?H?_?v?�?�?�?�?�? � �   00.0E0\0s0�0�0�0�0�0�01+1B1Y1p1�1�1�1�1�1�12(2?2V2m2�2�2�2�2�2�23%3<3S3j3�3�3�3�3�3�34"494P4g4~4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5686d6�6�67<7N7�788H8q8�8�8�8�8�89@9t9�9�9:2:�:�:�:�:;.;L;�;�;7<E<q<�<�<�<�<�<�<=&=4=I=]=o=�=�=�=�=�=�=�=>&>8>I>Z>k>|>�>�>�>B?l?�?   �   $0D0�0�0d1h1l1p1t1�12*2A2_2�2�2�3�3�3�3G4�45 5<5G5`5v5�5�5�5�5�5�56!6,6E6[6q6|6�6�6�6�6 787@7N7g7r7�7�7�78838|8�8�89 9<9R9c9o9}9�9�9�9�9:N:v:�:�:�:	;;5;K;a;�;�;�;<<(<n<}<�<�<�<�<�<�<=-=7=Q=p=�=�=�=�=�=>>>M>l>�>�>�>�>�>�>�>?>?M?W?q?�?�?�?�?�?�? � L  0N0]0|0�0�0�0�01-181Q1g1r1�1�1�1�12!2N2]2y2�2�2�2�2�233+363O3n3y3�3�3�3�3�3�34-474Q4g4�4�4�4�455%505I5Z5f5t5�5�5�5�56%6;6Q6g6}6�6�6�6�67 7<7G7`7q7}7�7�7�7�7�7818Q8o8�8�8�8�8�8�819@9\9r9�9�9�9�9�9�9:5:?:J:d:�:�:�:�:;;/;E;x;�;�;�;<<1<G<~<�<�<�<�<�<=!=,=E=d=z=�=�=�=�=�=	>>2>l>}>�>�>�>�>?-?L?W?p?{?�?�?�?�?   � �   0090O0e0{0�0�0�0�0�0�01+1A1W1m1�1�1�1�1�1�12232I2_2u2�2�2�2�2�2�23%3;3Q3g3}3�3�3�3�3�344-4C4Y4o4�4�4�4�4�4�4	5555K5a5w5�5�5�5�5�5�56'6=6S6i66�6�6�6�6�677/7E7[7q7�7�7�709e:�:�:�:�:�:�:�:�:;);~;�;�;�;A<c<�<�<	=�= >�>w?�?�?   � �   !070�0�0�01@1d1�1�1%2I2u2�2�2�2�23333Q3�3�3�3�3�3�3!424>4L4]4�4�4�4�4�455*5m5�5�5�5�5$6`6{67.7S7m7�7�78B8Z8v8t9�9�9�9Z:�:�:�:�:;;F;�;�;�;�;�;\<�<�<
=='=5=F=x=�=�=(>]>n>z>�>�>�>?)?4?[?f?�?   � �   0�0 1-1F1_1i1�1�1�1�1�1�1	2(2>2Z2p2�2�2�2�2�2�2
3)333O3
5O5;6�7�7�7�7�7�7�7�7 888|8�89y9�9�9�:;�;�;�;�;<,<8<F<�<�<�<�<�<�<�<
=V=�=
?\?|?   � �   00A0{0�0�1�1�3�307P7w7�7�7�7�78848W8�8�8�8�8F9�9�9�9:':;:J:X:l:�:�:�:�:�:V;n;<&<S<g<v<�<�<�<�<�<=i=}=�=�=�=�=�=�=>A>R>^>l>�>�>�>�>�>?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�? � �   0000000020<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3�3�3�3�3�344404<4_4l4�4�4�4�4�4�45,5H5Y5j5{5�5�5�5�566$626C6O6r66�6�6�6�6�6�6+7?7[7l7}7�7�7�7�788%818?8P8\88�8�8�8�8�8�8989L9h9y9�9�9�9�9�9:$:5:A:O:`:l:�:�:�:�:�:�:;;H;\;x;�;�;�;�;�;<+<4<E<Q<_<p<|<�<�<�<�<�<�<=(=X=l=�=�=�=�=�=>>;>D>U>a>o>�>�>�>�>�>�>�>?'?8?h?|?�?�?�?�?   �  00,0K0T0e0q00�0�0�0�0�0�01171H1x1�1�1�1�1�12(2<2[2d2u2�2�2�2�2�2�2�233/3G3X3�3�3�3�3�3�3$484L4n4w4�4�4�4�4�4�4�45515B5Z5k5�5�5�5�5�5�546H6\6{6�6�6�6�6�6�6�6�67%7>7O7g7x7�7�7�7�7�78D8X8l8�8�8�8�8�8�8�8�89!959N9_9w9�9�9�9�9�9
::T:h:|:�:�:�:�:�:�:�:;;4;H;a;r;�;�;�;�;�;<<.<d<x<�<�<�<�<�<�<�<�<=,=A=U=n==�=�=�=�=>>*>;>�>�>�>�>�>�>�>???B?O?d?x?�?�?�?�?�?    �  0+0<0M0^0�0�0�0�0�0�011#1/1R1_1t1�1�1�1�1�122;2L2]2n2�2�2�2�2�233"333?3b3o3�3�3�3�3�3�34/4K4\4m4~4�4�4�4�455$525C5O5r55�5�5�5�5�5�5+6?6[6l6}6�6�6�6�677'737A7R7^7l7}7�7�7�7�7�7�7�78'8t8�8�8�8�8�899+9M9V9g9s9�9�9�9�9�9�9�9�9 ::-:>:S:g:�:�:�:�:�:	;C;W;k;�;�;�;�;�;�;�;�;�;	<<(<@<T<m<~<�<�<�<=='=8=I=�=�=�=�=�=�=�=>>>,>=>I>W>h>�>�>�>�>�>�>4?E?V?g?x?�?�?�?�?   �  00'030A0R0^0l0}0�0�0�0�0�0�0�01'1t1�1�1�1�1�122+2M2V2g2s2�2�2�2�2�2�2�2�2 33-3>3S3g3�3�3�3�3�3	4C4W4k4�4�4�4�4�4�4�4�4�4	55(5@5T5m5~5�5�5�566'686I6�6�6�6�6�6�6�6777,7=7I7W7h7�7�7�7�7�7�748E8V8g8x8�8�8�8�899'939A9R9^9l9}9�9�9�9�9�9�9�9:':t:�:�:�:�:�:;;+;M;V;g;s;�;�;�;�;�;�;�;�; <<-<><S<g<�<�<�<�<�<	=C=W=k=�=�=�=�=�=�=�=�=�=	>>(>@>T>m>~>�>�>�>??'?8?I?�?�?�?�?�?�?�?   0 �  000,0=0I0W0h0�0�0�0�0�0�041E1V1g1x1�1�1�1�122'232A2R2^2l2}2�2�2�2�2�2�2�23'3t3�3�3�3�3�344+4M4V4g4s4�4�4�4�4�4�4�4�4 55-5>5S5g5�5�5�5�5�5	6C6W6k6�6�6�6�6�6�6�6�6�6	77(7@7T7m7~7�7�7�788'888I8�8�8�8�8�8�8�8999,9=9I9W9h9�9�9�9�9�9�94:E:V:g:x:�:�:�:�:;;';3;A;R;^;l;};�;�;�;�;�;�;�;<'<t<�<�<�<�<�<==+=M=V=g=s=�=�=�=�=�=�=�=�= >>->>>S>g>�>�>�>�>�>	?S?g?{?�?�?�?�?�?�?�?�?   @ �  00'080P0d0}0�0�0�011&171H1Y1�1�1�1�1�1�122"2.2<2M2Y2g2x2�2�2�2�2�2�2D3U3f3w3�3�3�3�3�34&474C4Q4b4n4|4�4�4�4�4�4�4�45#575�5�5�5�5�5�56'6;6]6f6w6�6�6�6�6�6�6�6�6�67$7=7N7c7w7�7�7�7�788S8g8{8�8�8�8�8�8�8�8�899'989P9d9}9�9�9�9::&:7:H:Y:�:�:�:�:�:�:;;";.;<;M;Y;g;x;�;�;�;�;�;�;D<U<f<w<�<�<�<�<�<=&=7=C=Q=b=n=|=�=�=�=�=�=�=�=>#>7>�>�>�>�>�>�>?'?;?]?f?w?�?�?�?�?�?�?�?�?�?   P �  0$0=0N0c0w0�0�0�0�011S1g1{1�1�1�1�1�1�1�1�122'282P2d2}2�2�2�233&373H3Y3�3�3�3�3�3�344"4.4<4M4Y4g4x4�4�4�4�4�4�4D5U5f5w5�5�5�5�5�56&676C6Q6b6n6|6�6�6�6�6�6�6�67#777�7�7�7�7�7�78'8;8]8f8w8�8�8�8�8�8�8�8�8�89$9=9N9c9w9�9�9�9�9::S:g:{:�:�:�:�:�:�:�:�:;;';8;P;d;};�;�;�;<<&<7<H<Y<�<�<�<�<�<�<=="=.=<=M=Y=g=x=�=�=�=�=�=�=D>U>f>w>�>�>�>�>?-?6?G?S?a?r?~?�?�?�?�?�?�?�?   ` |  0030G0�0�0�0�0�0�0#171K1m1v1�1�1�1�1�1�1�1�1�12 242M2^2s2�2�2�2�233)3c3w3�3�3�3�3�3�3�3�344)474H4`4t4�4�4�4�45%565G5X5i5�5�5�5�5�566!626>6L6]6i6w6�6�6�6�6�6�67T7e7v7�7�7�7�7�78-868G8S8a8r8~8�8�8�8�8�8�8�89939G9�9�9�9�9�9�9#:7:K:m:v:�:�:�:�:�:�:�:�:�:; ;4;M;^;s;�;�;�;�;<<)<T<i<u<�<�<�<�<�<=&=D=Y=e=u=�=�=�=�=>>4>I>U>e>�>�>�>�>�>?$?9?E?U?t?�?�?�?�?�?   p �   0)050E0d0t0�0�0�0�011%151T1d1u1�1�1�1�1	22%2D2T2e2q2�2�2�2�23373G3X3d3�3�3�3�34474G4X4d4�4�4�4�45575G5X5d5�5�5�56>6�6�6�6�6	7C7�7�7�7�7=8e8t8�8w:�:�:�:�:�:	;�;�;D<r<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=�=J>j>�>�>�> � �  1z1�1�1�1�1�1�1222B2g2t2�2�2�2�2�23)393^3n3�3�3�3�3�3424B4g4t4�4�4�4�4�45 5-5L5\5�5�5�5�5�5�5 606U6e6�6�6�6�6�67)797[7k7�7�7�7�7�7888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8 999?9S9e9y9�9�9�9�9�9::.:\:v:�:�:�:�:;;/;C;Q;�;�;�;�;�;<<<A<N<m<z<�<�<�<�<�<�<='=C=S=q=�=�=�=�=�=�=�=�=�=�=�=&>7>C>Q>r>y>�>�>�>�>�>�>?#?0?L?Y?q?�?�?�?�?�?�?�?�?�?   �   0+070E0W0j0~0�0�0�0�0�0�011/1d1�1�1�1p3�34;4^4�4�45555E5X5d5r5�5�5�5�5�5�5�5�56*6Q6e6w6�6�6�6�6�67&7B7]7q7�7�7�7�7�7�7818B8S8�8�8�8�8�89"9C9T9`9n9�9�9�9�9�9�9�9:j:{:�:�:�:�:�:�:�:6;G;S;a;�;<<I<c<�<�<,=�=�=�=�=�=g>�>�>�>�>�>�>??-?9?G?m?�?�?�?�?�?�?   � �   0!030G0`0{0�0�01�12F2f2�2�2�2�3�34�4	5-5A5h5�5�5y6�6�6�6�6�67_7r7�7�7�7�7�8�859�9t:�:�;�;�;
<</<@<m<�<�<�<�<�< ===/=C=U=f=w=�=�=�=�=�=�=>>/>@>Q>b>�>�>�>�>�>??=?Q?c?�?�?�?�?�?�?�?   �   0"030D0Y0m0�0�0�0�0�0�0�011/1g1v1�1�1�1�1 2 2+2J2h2�2�2�2�23)3M3�3�3�3�3�3�3H4Y4�4�4�4g5v5�5�56/6Q6�6�6�6�67.7J7�7�7�7�78808;8Z8x8�8�89W9f9p9�9�9�9�9�98:G:Q:q:�:�:7;F;k;�;�;�;�;�;�;<<W<f<p<�<�<�<�<==:=_=�=�=�= >%>D>f>�>�>�>�>�>?G?V?`?�?�?�?�? � �   030U0`00�0�0�0�0�01(1G1R1q1|1�1�1�12202\2�2�2�2�2	3333�3�3�3�344!4A4f4�4�4�4�455:5�5�5�5�56(6M6X6w6�6�6�6�67@7|7�7�7�78878U8�8�8�8�8�89q9�9�9�9:6:w:�:�:�:�:�:�:;9;�;�;�;<H<W<o<�<�<�<*=O=l=�=�=�=�=�=
>>4>?>�>�> � �   �0�0%1{1�1�12)2a2_6�6�8�8�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :b:�:�:;;P;�;<6>F>�>g?�?   � |   �0�0�0�0�0�0�0�0$1<1�1�1�12%2\3`3d3h3�3>4�4�455h5l5p5t5x5|5�5�7�7�8�8 9�9�:$;;;z;<p<t<x<|<�<�<�<6=G>i>�>�>?5?R? � t   �0�0�0�0�0�01�1282}2g344<4l4,5�56F6r6�6�6�6�6=7�7:8�8�9�9�9�9�9�9�9�9�9�:4;�;�;�<^=�=>Q>�>�>?.?`?h?�?     �   80<1@1D1H1�2�2�2I3U3h3�3�3�3\4h4{4�4�4�425>5Q5�6�6~7�7888@8p8�9�9�9�9�9:X:�:�:�:�:8;t;|;�;�;�;�;T<=�=�=�=�=�=8>�>�>�>?s?�?    �   0!0O0�0�0"1R1~1�1�1;3�3t4x4|4�45U5�57768�8�8�8�8�879?9�9�9�9:8:�;�<|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>'>r>�>�>�>�>?&?�?�?�?�?     |   R0j0�0 101\1|1�1�1`4d4h4l4p4t4x4|4�4�4�45L5x5�5�5�5�56�6�6778�8�8�8�89�9�9�9�:�:;_;j;�;�;<><�<�<�<?=v=�=0>? 0 l   C2T2m2�2�2'3�3d4�4T5�6�6r7�9�9�9K:�:�;�;<D<t<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<D=N=e=�=>Q>~>�>�? @ �   1�1�23'4W4�4�4�4E5�56666[6�6�78+8C8[8�8�8�89#9G9Z9f9t9�9�9�9�9�9::0:B:S:h:�:�:�:�:�:;&;:;L;];r;�;�;�;�;�;<�<�<�<==d=�=�=�=�=>>A>f>�>�>�>�>�>'?6?�?�? P   0040H0\00�0�0�0�0�01/1C1R1d1�1�1�1�1�12#222D2q2�2�2�2*3G3g3�3�3�3�34.4w4�4�4�45#5T5f5�5�5�56#6a6u6�6�67D7t7�7�7�7�7�7�7�7�78838D8U8f8x8�8�8�89.9=9U9o9�9�9�9:H:q:�:�:�:�:�:';:;d;s;�;�;�;�;�;�;<)<?<P<\<j<�<�<�<=g=�=�=�= >>1>B>N>\>z>�>�>�>�>?:?]?n?z?�?�?�?   `   0$0?0u0�0�0�0�051d1s1�1�1�12"2H2^2|2�2�2�2�23$3@3Z3�3�3�3�3�3@4O4q4�4�4�4�4�4D5[5l5~5�5�5�5�5�5�5
66(606D6H6L6P6T67.7=7c7�78~8�89*9o9�9�9�9�:�:�: ;;A;[;w;�;�;�;�;�;�;<4<N<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<N=~=�=�=�=�=>5>M>`>�>�>�>�>�>?%?=?P?s?�?�?�?�?�? p   0-0@0c0{0�0�0�0�0�0101S1k1~1�1�1�1�12+2>2N2c2{2�2�2�2�2�2�23.3F3Y3�3�3�3�3�3�34(4>4N4c4{4�4�4�4�4�4�45535K5`5v5�5�5�5�5�5�566D6u6�6�6!717A7Q7w7�7�7�7Q8`8j8�8�899t9�9�9�9':>:�:�:�:�:;.;w;�;�;�;�;&<1<d<x<�<�<�<=9=g=x=�=�=�=>">�>�>Y?m?�?�?�?�?�? �   0+0D0X0q0�0�0�0�0�01 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1�12C2d2�2�2�2�2�2 3#3A3T3w3�3�3�3�3�34+4>4a4y4�4�4�4�455.5Q5i5|5�5�5�5�566A6_6r6�6�6�6�6�67707F7V7k7�7�7�7�7�7�7%8K8`8v8�8�8�8�8�8�89909F9V9k9�9�9�9�9�9�9 ::&:;:S:h:~:�:�:�:8;�>�>�>�> � �   �2�2�2�2	3&3<3�3�3�3�34G4j4�4�4�4�4�4�4�5�5�5�5�56C6x6�6�6�6�6,7074787<7@7D7�7�78"8R8q8�8�8�899$9a9t9�9�9�9�9:!:4:T:|:�:+;L;f;�;�;�;�;4<Q<�<�<=$=Q=b=�=�=�=�=�=�=>>#>A>R>t>�>�>�>�> ??4?T?l?�?�?�?�?�?�?   �    000/0c0v0�0�0�0�0�0�01$1D1d1�1�1�1�1�1$262D2V2t2�2�2�2�23 3D3a3t3�3�3�3�34!414D4d4�4�4�4�45$5D5d5�5�5�5�56W6�6�6�6�6�6-7d7}7�7�7�7�7$8B8]8t8�8�8�89-9D9[9r9�9�9:$:D:d:�:�:�:�:;0;D;V;v;�;�;�;�;�;0<D<�<�<�<=(=H=�=�=�=�=>*>�>�>�>�>?4?�?�?�?�? � $  0$0T0q0�0�0�0�0�0�0�011-1<1N1q1�1�1�1�1�122,2>2d2~2�2�2�2�23$3D3d3�3�3�3�34$4D4d4�4�4�45$5D5d5�5�5�5�56$6D6d6�6�6�6�6747T7t7�7�7�7�7848T8t8�8�8�8�8949T9t9�9�9�9�9:;:d:�:�:�:�:�:;1;D;a;q;�;�;�;�;�;�;<$<D<d<�<�<�<�<=6=N=x=�=�=�=�=>$>D>d>�>�>�>�>�>�>�>$?>?R?`?o?�?�?�?   �    00+090P0d0}0�0�0�0�0�01141T1t1�1�1�1�12$2A2d2�2�2�2�23$3D3d3u3�3�3�3�34T4�4�4�4�45$5A5T5t5�5�5�5�56>6�6�6�6�67D7a7�7�7�7�7�78$8D8d8�8�8�8�8�8�89949T9t9�9�9�9�9!:4:T:t:�:�:�:�:;E;Z;k;�;�;�;�;C=J=Q=X=_=f=m=t={=�=�=�=�=�=�=�=�=X>i>u>�>   � �   00$0+02090�0�0�0�01R1t1�1�1�1222F2V2�2�2�2�233!313A3T3�3�3�3444Q4d4�4�4�4�45D5g5�5�566+6g6�6�6�6�6747T7q7�7�7�7	818D8w8�8�8�8 9�9�9�9:t:�:�:�:�:�:(<S<�<==�=�>?1?D?a?t?   � �   �1�1�1�1�2�24�4�4$5*505<5A5f5m5�5�5�5*686o6�6�6�6�6�6�6S7m7�7�7�78!848Q8d8�8�8�8�8 9t9�9:�:�:�:�:;�;<'<p<�<�<�<=1=Q=t=�=�=�=>$>D>d>�>�>�>�>�>?4?T?t?�?�?�?�?�?   � �   "060J0f0~0�0�0�0�01111=1g1�1�1�12G2�2�23T3t3�3�3�3474a4�4�4�4545T5�5�5�56*6W6�6�6�6777i7�7�7�7<8w8�8�8�8�8�89!9�9�91:;-;k;�;�;�;
<4<Q<q<�<�<�<7=d=�=�=�=h>�>�>�>�>�>?&?O?a?�?�?�?   �   0%0G0�0�0�0�0�0�1�1�1�1:2�2�2@3`3�34454L4b4�4�4�4�45B5T5�5�5;6�6�6737b7�7�78K8�8�8�8�8$9_9�9�9:W:�:g;�;�;�;�;7<^<�<�<4=L=n=�=�=�=�=>K>�>�>�>)?v?�?�?�?    �   '0A0y0�0�01?1Z1�1�1�12:2\2p2�2�23�4�4�4�4,56-6L6i6�6�6�617q7�7�78'8T8�8�8�89d9�9:d:�:;T;�;�;D<�<�<4=�=�=$>q>�>?T?�?�?     �   ;0�0�0	1t1�1�1!2k2�2�23D3{3�3�3444~4�45a5�5�5�5�56G6w6�6�6/7o7�7�7-8d8�8�8�89D9t9�9�9:Q:�:�:�:!;Q;�;�;�;�;q<�<�<�<=2=q=�=�=�=�=>/>A>�>�>�>�>?? ?<?X?a?�?�? 0 �   '0D0y0�0u1�1H2L2P2T2X2\2`2d2h2�2b3�3�3�3�3�3�3�3�3�3�4�4�4�4�4�45X5�5�5�5�5�56D6p687W7A8�89f9�9�9�9:$:D:X:h:�:�:�:�:;; ;7;L;`;};�;�;�;�;�;�;<D<d<�<�< =%=6=Q=w=�=�=�=>>B>]>p>�>�>�>?r?�?�?�?�? @ �   00(0>0C0h0|0�0�0�0�0�011'1H1\1�1�1�1�1242�2�2�23E3�3!4&4B4^4t4y4�4�4�4�45C5�5�5�5@6^6�6�6�6�6737E7V7k7|7�7�7�7�78;8q8�8�8�839Q9�97:U:�:�:�;�;W<^<�<=%=>#>k>t>�?   P �   000T0t0�0�0�01$1A1a1�1�1�1�1~2�2�2�23$3Q3�3�3�34)4H4�4�4�45^5j5�5�56696p67�7p8�8�89	99m99�9�9�9�9::d:�:�:�:�:5;Q;{;�;�;�;�;1<9<I<j<�<�<�<==9=�=�=�=
>>K>Y>q>�>�>�>�>�>�>�>???#?1?C?n?�?�?�? ` �   "0T0X0\0`0d0h0�0�0�0	11%1-171E1M1e1o1y1�1�1�1J2V2u2734�4�4�5�67�7�7`8d8h8l8p8t8G9�9�:�:�:;;�;"<J<}<�<�<v=�=">o>�>�>?'?B?�?�?�? p �   0*0�0�0�01k11�1�12�2�2�2�2�2�2�3-4S5]5�5�6I7�7V9^9�9�9�9�9�9�9�9:>:�:�:�:�:�:*;5;=;b;�;�;<3<�<�<=="=0=g=�=�=�=%>�>�>�>�>�>�>A?P?�?�?�?�? � �   00#0Z0b0�0�0�0�0�01'1T1�1�1�1�1�1?2M2�2�2�23D3d3�3�34G4w4�4�4545T5q5�5�5Z6�6�6�67J7t7�7�7�78#8�8�8�8
9;�;,<q<�<�<�<
=1=T=�=�=�=�=>D>d>�>�>�>�>?4?g?�?�?�?�?   � �   0D0d0�0�0�0�01$1D1d1�1�1�1�1�1242Q2t23*3�3&4G4�4�4'5�5�56�6�6E7�7�7a8�8�89)9g9�9M:i:�:�:�:<;d;�;=<Y<t<�<�<,=�=�=�=�=7>�> ?:?�? � �   -0I0d0y0�01�1�112�2�2D3�3�3�3�3414T4�4�4�4525e5�5�5�5�5�5!6A6d6�6�6�6�6�6!7A7g7�7�7�7$8A8T8t8�8�8�8�8919P9U9Z9_9t9�9�9�9�9:$:T:k:�:�:�:;';W;�;�;<G<<�<�<�<=q=�=�=�=�='>Q>d>�>�>�>?'?T?t?�?�?�? �   $0G0�0�0�0�0�0�01$1A1Q1d1�1�1�1�1242H2T2b2s2�2�2�2�2�2�2343N3b3r3�3�3�3�3�3444T4t4�4�4�4�45!515D5d5�5�5�5�5606T6t6�6�6�6�67$7D7�7�7�78$8D8d8�8�8�8�8�8949T9t9�9�9�9�9�9::4:T:w:�:�:4;T;t;�;�;�;�;<4<t<�<�<�<�<=!===I=�=�=>A>d>�>�>�>?$?T?�?�?�?�? �    080]0~0�0�0�01,1@1P1t1�1�1�12$2<2\2�2�2�2�233=3d3w3�3�3�3�3�3%4=4]4�4�4�4�4�45-5E5e5�5�5�5�56%6E6l66�6�6�67.7T7t7�7�7�7�78$8D8d8�8�8�8�8�8949T9t9�9�9�9�9:4:T:t:�:�:�:�:�:;4;T;t;�;�;�;<D<q<�<�<�<�<=1=T=t=�=�=�=>J>�>�>�>?1?W?�?�?�?   � �   0)0a0�0�0�0�0�081W1w1�1�1�1�12$2N2_2�2�2�2�2373a3�3�3�3�3414Q4t4�4�4�4$5T5�5�5�56$6Q6q6�6�6�6747d7�7�7�7�78A8a8�8�8�8�89G99�9�9::�:;?;S;l;�;�;�;<:<\<�<�<�<$=Q=q=�=�=�=�=>4>d>�>�>�>�>?4?R?p?�?�?�?   � �   !0D0q0�0�0�0�01141�1�1�1'2T2t2�2�213T3�3�3�3494P4n4�4�4�4�5�5�5 6;6@6g6�6�8�:�:=;J;~;�;�;�;<x=|=�=�=�=�=�=>D>d>�>�>�>�>?)?k?�?�?�? � �   0Y0�01D1�1�1�1�112T2q2�2K3P3Q6q6�6�6�6�6747W7�7�7�7�78$8D8{8�89W9�9�9D:�:�:�:�:�:�:�:;;�;�;�;�;�<=�=�=>>�>�>�>?!?G?w?�?�?�?     0  00$0-0>0h0m0�0�0�0!1G1t1�1�1�1�142�2�23�3�3464w4�4�4�45#5/5A5X5j5{5�5�5�5�5�56'686K6u6�6�6�6�6�6�6�6�67(7A7m7�7�7�7�7�7�78808C8e8t8�8�8�8�8�8�8�89919]9w9�9�9�9�9�9�9: :,:::\:m:�:�:�:�:�:;;";8;J;[;g;u;�;�;�;�;<<$<2<T<e<�<�<�<�<�<�<�<=7=H=T=b=�=�=�=�=�=�=>4>�>�>�>0???J?X?j?�?�?�?  �   0$060G0n0�0�011111�1�1�1�1�1�1212M2�2�2�2�2�2�233+3}4�4�4�4�4�4�4�4�4�4�4�5d6n6x6�6�6�6�6�6�6�6�8�8�8�8%9;9�9 :::::#:*:1:8:?:F:";U;y;�;�;5<Y<�<�<�<===e=�=�=�=5>r>�>�>�>%?e?�?�?   �   "0G0f0�0�0191a1�1�1�1�1�1292h2�2�23F3k3�3�3-4u4�4�4"5U5�5�56E6�6�67U7�7�7858u8�8�8B9u9�9�9:P:�:�:%;e;�;�;5<u<�<=8=S==�=�=�=�=">b>�>�>?�?�? 0 �   0H0�0�0�01H1�1�1�152r2�2�223r3�3�3$4r4�4�455t5q6�6�67X7�78E8�8�89E9�9�9:E:�:�:�:";R;�;�;%<e<�<�<5=�=5>�>�>?U?�?�?�?�?�?�?�?�? @ �   0U0�0�01R1�1�152u2�2d3�3�3�3474R4~4�4�45,5E5s5�5�5616d6�6�6�67J7�7�7*8?8~8�8�8�8J9m9�9�9�9�9�98:j:�:�:�:�:$;t;<2<h<�<�<�<�<=5=u=�=�=>U>�>�>%?e?�?   P �   0B0�0�01U1�1�12$21272h2�2�2�2�2 333333,343T3�3�3$4T4z4�4�4�4+575�5�5�566)6A6�6�6�6�6�6 77747\7o7t7�7�7�7�7�7Q8t8�8�8�89!9D9T9�9�9�9�9:$:Q:q:�:�:�:�:;4;T;�;�;�;�;<1<T<t<�<�<$=d=�=�=>$>D>d>�>�>�>�>?1?T?�?�?�? ` <   *0Q0t022G2L233M3R344F4K4�4�4X7�7�=>> >$>(>   p `   �0�0�0�01�3�6�6�6%7e7�7�7%8b8�8�89B9u9�9�95:r:�:�:;2;e;�;�;%<e<�<�<%=e=�=>U>�>�>%?u? � �   0,020�0�0�01.1�122l2y2�2�2�2�2�3�3�3�3�3�3W4c4k4w4�4�4�45575Y5�6�6�6�6"7*7>7H7f7r7~7�7�7�7�7�7�7�7	88!8N8X8`8�8�8�8�8�8�8�8�8979J9f9z9�9�9<:H:X:d:�:�:�:�:;;�;�;�;�;<F<R<s<�<�<=�=�='>3>b>�>�>�>??H?^?t?}?�?�?�?�?�?�?�?   � �   -0�0�0�0&121J1R1�1�12�2�2�2�2Q3Y33�3�3�3�3+4�4�4�4^5f5�5�5�5\6�6�6Z7n7�7�7�7�79;9C9P9<:H:X:d:�:�:�:�:;;~;�;�;�<
=#=�=�=�=�=�=*>C>�>�>�>�>3?[?i? � (  131L1S1[1`1d1h1�1�1�1�1�1�1�1�1�1�1�1B2H2L2P2T2�2�2�2�2�2�2�23?3q3x3|3�3�3�3�3�3�3�3�3�3�3�3t5�5�556;6?6D6J6N6T6X6^6b6g6m6q6w6{6�6�6�6�6�6�6�6�67'717;7|7�7�7�7,8A8[8�8�8l9r9�9�9�9�9�9S:{:�:5<S<l<s<{<�<�<�<�<�<�<�< =======b=h=l=p=t=�=�= >>>>>5>_>�>�>�>�>�>�>�>�>�>�>????   � �   �0�0�0�0�0L1Y1�1�1�12!2`2l2�2�2�2�23#3+3�3�3�3�344#4X4a5i5q5A6I6Q6Y6w66�6�6777�7�7�7�7�7�7�8�8�8�8�89
9z99�9�9�9�9�9�9):9:;[;f;l;�<�<?=F=\=f=�=S>Z>�>�>�>?3? � �   �2n3�4�4553595�6�899
99999:H:\:�:�:�:�:�:�:�:�:;;;;;#;*;1;8;@;H;P;\;e;j;p;z;�;�;�;�;�;�;!<�<*=:=F=X=h=t=y>�>�?�?   � �   0-0D0O0~0�0�0�01-1B1L1e1o1|1�1�1�1�1�1%2c2�2�2�2�2�2�2	33!373b3|3�3�3�3�3�3�3�3�3�3�3 4C4G4K4O4S4W4[4_4c4g4k4o4s4w4�4�4E5W5�5�5�5�56y6�6�6�6�6�6�627�7�7�7�7�7�78"8^8�8�8�8�8�9�9�9�9�:;";B;�;�;�;	<<A<L<^<�<�<===2=H=�=>�>   � D   ?0`0e0�5�5&6�7�8w;};�;=�=�=�=�=C>]>�>�>�>�>�>�>?3?u?�?�?�? � �  0&070K0S0\0e0�0�0�0�0�0�0�0�0�0�0111)191>1C1T1Y1j1o1|1�1�1�1�1�1�1�1222 2*2@2a233%313A3G3X3w3�3�3�3�3�3�3�3�3 4/464D4M4�4�4�4�4�45>5s5�5�5�5�556m6�6�67!7G7W7l7v7|7�7�7�7�7�9�9�9�9:#:/:>:I:o:�:�:�:�:�:�:�:;7;];q;|;�;�;�;�;�;�;�;�;�;�;�;<<<,<<<E<M<e<x<~<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<=====$=,=1=7=?=D=J=R=W=]=e=j=p=x=}=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>#>(>.>6>;>A>I>N>T>\>a>g>o>t>z>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>???*?3?X?m?�?�?�?   �    00070<0a0~0�0k1s1�1�1�1Y2_2�2�2�2�2�2-3E3O3k3r3x3�3�3�3�3�3�3�3�3�3424�4 5b5�5#656[6~6�6�6�6�6]7w7�7�7�7�7�7�8�8�8 99999$9w9|9�9�9�9�9�9�9�9F:P:k:u:�:P;y;�;�;�;�;h<o<�<�<�<�<�<�<�<�<�<=	== =F=w=�=�=�=�=&>:>_>�>�>�>Y?�?  �   M0�0�0�0$1�1 2)22�2e3p3�3�3Y4b4n5w5c6�6�6�687o7�7�78+8�8�8
9$9�9:�:�:�;�;<F<�<�<�<�<=
==)=8=B=O=Y=i=�=�=	>y?�?�?�?�?�?   �   0�0�0�0�0�01-1H1P1^1c1r1�1�1282K2�2363�3�4�4x5�5�6Q7�7�7�78!8M8U8x8�8D9\9p9�9�9�9:%:-:9:�:�:�:�:�:;(;t<|<�<�<{=|>�>�>�>�>�>�>?? ?>?J?V?b?�?�?�?�?�?�?�?�?   0 �    040>0F0g0{0�0�0�0�0�0�0�0$131;1A1X1^1o1�1�1�122!2>2D2Y2~2�2�2N3�3�3�3�3�3�34?4K4�4�5�5�5�56�6�67H7e7y7�7�7S8[8�8�8�8�8�8999#9A9M9c9l9u9�9$:^:r:�:�:�:�:;4;�;N<_<�<�<�<�<$=H=Q=\=�=�=+>k>r>�>�>?i?�?   @ d   0G0�0�01141w1�2�2�2�2�3(4z4�4�45i5u5�5�5�5�5�5�536?6�6�6�6Z7�7�8�8�8�8�8�9�<w=�=f?q?�?�? P l   $060H0�0�0�0	1121H1Q1]1h1�1�1�12202E2K2u2�2�3	44w5�5�728�9�;�;<+<?<E<�<==!=-=�=�=�=%>=>�>�>�> ` �   }0�0�0�0�0�0�0�0111(1/1?1E1K1S1Y1_1g1m1s1{1�1�1�1�1�1�1�1�1�1�1�132K2d2�2�2�2$313]3e3�3�34E4Q4q4�4�4�4	555�5�5�5�566"6W6�7�7�7I8Q8Y8a88�8�8�8	99!9x9�9�9�9�9�9�9�:�:�:�:;;;�;%<0<R<�<�<�<I=U=|=�=�=�=�=>.>r>{>?K?�?�?�?   p h   010C0U0g0y0�0�0�0�0�0�0�01(1:1L1^1�4Y5�5�6=7z7�789�9�9::(:�:;;;+;Q;�;�<�<�>,?8?�?�?�?�? � T   u0�0�0:1\2d24�4�485@5L5[5�5�586�6 :2:�=�=�=�=�=�=�=�=�=�=�=�=�=�>�>�>�>?|? � $   �9[<�<====R=\=�=�=�=�=�=�? � (   00D0�0�01$1�1�1�1�1�1�122   � �  �011111$1(1,1x2|2�2�2�2�2�2�2�2�2D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444444l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555555 5$5(5,5054585<5@5D5H5L5P5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � x   00000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< � 0  h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3444444 4$4(4,4<4@4D4H4L4P4T4X4\4`4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5$5(5,5054585<5@5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$686<6@6D6H6L6P6T6X6\6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7$7(7,7074787�7�7�7�7�7�7�7�7�7�78888888 8$8(8@8D8H8L8P8T8X8\8`8d8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999$9(9,9094989<9@9D9H9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::::: :$:(:@:D:H:L:P:T:X:\:`:d:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;0;4;8;<;@;D;H;L;P;T;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<< <$<(<,<0<4<8<<<P<T<X<\<`<d<h<l<p<t<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=<=@=D=H=L=P=T=X=\=`=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>(>,>0>4>8><>@>D>H>L>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>??? ?$?(?,?0?4?8?P?T?X?\?`?d?h?l?p?t?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � �   00000000 080<0@0D0H0L0P0T0X0\0�0�0�0�0�0�0�0�0�0�0P1T1X1\1`1d1h1l1p1t1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222222 2$2(2@2D2H2L2P2T2X2\2`2d2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333333034383<3@3D3H3L3P3T3�3�3�3�3�3�3�3�3�3�3�3�3�5�5�5�5 6666666P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8   � (  �0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111122�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�6�6�6 7$7(7,70747�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9 `     3$3(3   �    �4�4 � L  |1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,2�;�;�;�; <<<<<<<< <$<(<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � �  0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888 8(80888@8H8P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h: �    D=H=L=P= �    j8n8r8v8 0 �   �:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<   ` �   l<p<�<�<�<�<==,=<=@=T=X=\=d=|=�=�=�=�=�=�=�=�=�=�=�=�=>>>> >(>@>D>\>l>p>t>x>�>�>�>�>�>�>�>�>�>�>�>????4?8?P?`?d?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   p l  00 0004080<0@0H0`0d0|0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111 1(1@1P1T1d1h1l1p1t1|1�1�1�1�1�1�1�1�1�1�1�12222 24282H2L2P2T2X2`2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33 30343D3H3L3P3T3\3t3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�344,404@4D4H4L4P4X4p4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55(5,5<5@5D5H5L5T5l5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56$6(686<6@6D6H6P6h6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67 7$74787<7@7D7L7d7t7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�788 8084888<8@8H8`8p8t8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8999,9094989<9D9\9l9p9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:::(:,:0:4:8:@:X:h:l:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;$;(;,;0;4;<;T;d;h;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<< <$<(<,<0<8<P<`<d<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<=== =$=(=,=4=L=\=`=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=>>>> >$>,>D>T>X>h>l>p>t>|>�>�>�>�>�>�>�>�>�>�>�>?????4?D?H?X?\?`?d?l?�?�?�?�?�?�?�?�?�?�?�?�?�?   � @   000$04080H0L0P0T0\0t0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01$1(181<1@1D1L1d1t1x1�1�1�1�1�1�1�1�1�1�1�1�1�1222(2,20242<2T2d2h2x2|2�2�2�2�2�2�2�2�2�2�2�2�23333 3$3,3D3T3X3h3l3p3t3|3�3�3�3�3�3�3�3�3�3�3�34444444D4H4X4\4`4d4l4�4�4�4�4�4�4�4�4�4�4�4�4�4 555$54585H5L5P5T5\5t5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56$6(686<6@6D6L6d6t6x6�6�6�6�6�6�6�6�6�6�6�6�6�6777(7,70747<7T7d7h7x7|7�7�7�7�7�7�7�7�7�7�7�7�78888 8$8,8D8T8X8h8l8p8t8|8�8�8�8�8�8�8�8�8�8�8�89999949D9H9X9\9`9d9l9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::$:4:8:H:L:P:T:\:t:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;$;(;8;<;@;D;L;d;t;x;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<(<,<0<4<<<T<d<h<x<|<�<�<�<�<�<�<�<�<�<�<�<�<==== =$=,=D=T=X=h=l=p=t=|=�=�=�=�=�=�=�=�=�=�=�=>>>>>4>D>H>X>\>`>d>l>�>�>�>�>�>�>�>�>�>�>�>�>�> ???$?4?8?<?@?H?`?p?t?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � �  000,0004080<0D0\0l0p0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111(1,1014181@1X1h1l1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 222$2(2,20242<2T2d2h2x2|2�2�2�2�2�2�2�2�2�2�2�2�23333 3(3@3P3T3d3h3l3p3x3�3�3�3�3�3�3�3�3�3�3 44444,4<4@4P4T4X4`4x4|4�4�4�4�4�4�4�4�4�4�4�4 555$5(585<5L5P5`5d5t5x5�5�5�5�5�5�5�5�5�5�5�5�5 66 60646D6H6P6h6x6|6�6�6�6�6�6�6�6�6�6�6�6�67X7t7x7�7�7�7�7 88(8H8h8�8�8�8�89$9(9H9d9h9�9�9�9�9�9�9:0:P:p: � P  $0(02222 2$2(2,20242�2�2T9X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<$<D<P<T<X<\<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=�>�>�>�>�>�>�>�>�>�>�>?????? ?$?,?0?P? � �   X2p2�2�2�2�2�23,3D3`3|3�3�3�3�34(4D4`4|4�4�4�4�45(5D5`5|5�5�5�5�5606L6h6�6�6�6�6�6787X7t7�7�7�7�78 8@8`8�8�8�8�8 9 9D9h9�9�9�9�9:<:\:|:�:�:�:;@;h;�;�;�;<@<h<�<�<�<=<=l=�=�=�=>H>t>�>�>�> ?L?x?�?�?   � H   0,0X0�0�0�0101X1�1�1�1242`2�2�2�23<3`3�3�3�3�34,4H4d4|4�4�4                                                                            